
module Adder_cntrl ( CLK, Datain1, Datain2, Data_valid, Dataout, Exc, Mode, 
        Debug, Adder_datain1, Adder_datain2, Adder_valid, Adder_dataout, 
        Adder_carryout, Adder_ack, ExcCheck_valid, Exc_value, Exc_Ack, 
        RSTn_BAR, Dataout_valid_BAR, ExcCheck_Datain_15_, ExcCheck_Datain_14_, 
        ExcCheck_Datain_13__BAR, ExcCheck_Datain_12_, ExcCheck_Datain_11_, 
        ExcCheck_Datain_9_, ExcCheck_Datain_8_, ExcCheck_Datain_6_, 
        ExcCheck_Datain_5_, ExcCheck_Datain_4_, ExcCheck_Datain_3_, 
        ExcCheck_Datain_2_, ExcCheck_Datain_1_, ExcCheck_Datain_0_, 
        ExcCheck_Datain_10__BAR, ExcCheck_Datain_7__BAR );
  input [15:0] Datain1;
  input [15:0] Datain2;
  output [15:0] Dataout;
  output [2:0] Exc;
  input [2:0] Mode;
  output [4:0] Debug;
  output [8:0] Adder_datain1;
  output [8:0] Adder_datain2;
  input [8:0] Adder_dataout;
  input [2:0] Exc_value;
  input CLK, Data_valid, Adder_carryout, Adder_ack, Exc_Ack, RSTn_BAR;
  output Adder_valid, ExcCheck_valid, Dataout_valid_BAR, ExcCheck_Datain_15_,
         ExcCheck_Datain_14_, ExcCheck_Datain_13__BAR, ExcCheck_Datain_12_,
         ExcCheck_Datain_11_, ExcCheck_Datain_9_, ExcCheck_Datain_8_,
         ExcCheck_Datain_6_, ExcCheck_Datain_5_, ExcCheck_Datain_4_,
         ExcCheck_Datain_3_, ExcCheck_Datain_2_, ExcCheck_Datain_1_,
         ExcCheck_Datain_0_, ExcCheck_Datain_10__BAR, ExcCheck_Datain_7__BAR;
  wire   N144, N145, N146, N147, N148, N149, N151, N152, N153, N154, N155,
         N156, N157, N158, N160, N161, N162, N164, N165, N166, Debug_valid_reg,
         Op1_Sign_reg, Op2_Sign_reg, Op2_Mantissa_reg_7_, exc_reg_0_,
         carry_reg, N252, N253, N254, N255, N256, N257, N258, N259, N270, N362,
         N363, N364, N365, N366, N368, N369, N418, N419, N420, N422, N424,
         N425, N691, N2921, N2923, n73, n103, n109, n110, n111, n112, n113,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n212, n213,
         n214, n215, n216, n217, n218, n219, n222, n223, n274, n277, n664,
         n672, n915, n922, n991, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1103, add_x_35_A_9_,
         add_x_35_A_8_, add_x_35_A_7_, add_x_35_A_6_, add_x_35_A_5_,
         add_x_35_A_4_, add_x_35_A_3_, add_x_35_A_2_, add_x_35_A_1_,
         add_x_35_A_0_, C1_DATA1_7, C1_DATA1_5, C1_DATA1_4, C1_DATA1_3,
         C1_DATA1_2, C1_DATA2_7, C1_DATA2_5, C1_DATA2_4, C1_DATA2_3,
         C1_DATA2_2, C1_DATA3_7, C1_DATA3_6, C1_DATA3_5, C1_DATA3_3,
         C1_DATA3_2, C1_DATA3_1, C1_DATA4_7, C1_DATA4_6, C1_DATA4_5,
         C1_DATA4_3, C1_DATA5_7, C1_DATA5_6, C1_DATA5_5, C1_DATA5_3,
         C1_DATA5_2, C1_DATA5_1, C1_DATA6_7, C1_DATA6_5, C1_DATA6_4,
         C1_DATA6_3, C1_DATA6_2, C1_DATA7_7, C1_DATA7_6, C1_DATA7_2,
         C1_DATA7_1, C1_DATA8_7, C1_DATA8_6, C1_DATA8_5, C1_DATA9_7,
         C1_DATA9_6, C1_DATA9_5, C1_DATA9_3, C1_DATA9_2, C1_DATA9_1,
         C1_DATA10_7, C1_DATA10_6, C1_DATA10_5, C1_DATA10_3, C1_DATA10_2,
         C1_DATA11_5, C1_DATA11_4, C1_DATA11_3, C1_DATA11_2, C1_DATA11_1,
         C1_DATA11_0, C1_DATA12_5, C1_DATA12_3, C1_DATA12_2, C1_DATA12_1,
         C1_DATA12_0, C1_DATA13_5, C1_DATA13_4, C1_DATA13_3, C1_DATA13_2,
         C1_DATA13_1, C1_DATA13_0, C1_DATA14_7, C1_DATA14_5, C1_DATA14_4,
         C1_DATA14_3, C1_DATA14_2, C1_DATA14_1, DP_OP_979_173_2805_n80,
         DP_OP_979_173_2805_n79, DP_OP_979_173_2805_n78,
         DP_OP_979_173_2805_n77, DP_OP_979_173_2805_n76,
         DP_OP_979_173_2805_n58, DP_OP_979_173_2805_n55,
         DP_OP_979_173_2805_n52, DP_OP_979_173_2805_n48,
         DP_OP_979_173_2805_n45, DP_OP_979_173_2805_n44,
         DP_OP_979_173_2805_n43, DP_OP_979_173_2805_n39,
         DP_OP_979_173_2805_n35, DP_OP_979_173_2805_n20,
         DP_OP_979_173_2805_n19, DP_OP_979_173_2805_n18,
         DP_OP_979_173_2805_n17, DP_OP_979_173_2805_n16,
         DP_OP_979_173_2805_n15, DP_OP_979_173_2805_n14,
         DP_OP_979_173_2805_n13, DP_OP_979_173_2805_n12,
         DP_OP_979_173_2805_n11, DP_OP_979_173_2805_n10, DP_OP_979_173_2805_n9,
         DP_OP_979_173_2805_n1, DP_OP_989_183_2805_n55, DP_OP_989_183_2805_n48,
         DP_OP_989_183_2805_n43, DP_OP_989_183_2805_n38,
         DP_OP_989_183_2805_n26, DP_OP_989_183_2805_n25,
         DP_OP_989_183_2805_n23, DP_OP_989_183_2805_n14,
         DP_OP_989_183_2805_n13, DP_OP_989_183_2805_n12,
         DP_OP_989_183_2805_n11, DP_OP_989_183_2805_n10, DP_OP_989_183_2805_n9,
         DP_OP_989_183_2805_n8, DP_OP_989_183_2805_n5, DP_OP_989_183_2805_n4,
         DP_OP_989_183_2805_n3, DP_OP_989_183_2805_n2, DP_OP_989_183_2805_n1,
         DP_OP_990_184_2805_n58, DP_OP_990_184_2805_n51,
         DP_OP_990_184_2805_n48, DP_OP_990_184_2805_n43,
         DP_OP_990_184_2805_n34, DP_OP_990_184_2805_n26,
         DP_OP_990_184_2805_n25, DP_OP_990_184_2805_n23,
         DP_OP_990_184_2805_n22, DP_OP_990_184_2805_n21,
         DP_OP_990_184_2805_n14, DP_OP_990_184_2805_n13,
         DP_OP_990_184_2805_n11, DP_OP_990_184_2805_n10, DP_OP_990_184_2805_n9,
         DP_OP_990_184_2805_n5, DP_OP_990_184_2805_n2, DP_OP_991_185_2805_n48,
         DP_OP_991_185_2805_n43, DP_OP_991_185_2805_n38,
         DP_OP_991_185_2805_n14, DP_OP_991_185_2805_n11,
         DP_OP_991_185_2805_n10, DP_OP_991_185_2805_n9, DP_OP_991_185_2805_n5,
         DP_OP_991_185_2805_n4, DP_OP_991_185_2805_n3, DP_OP_991_185_2805_n2,
         DP_OP_992_186_8739_n32, DP_OP_992_186_8739_n31,
         DP_OP_992_186_8739_n30, DP_OP_992_186_8739_n29,
         DP_OP_992_186_8739_n23, DP_OP_992_186_8739_n19,
         DP_OP_992_186_8739_n17, DP_OP_992_186_8739_n16,
         DP_OP_992_186_8739_n15, DP_OP_992_186_8739_n13,
         DP_OP_992_186_8739_n12, DP_OP_992_186_8739_n11, DP_OP_992_186_8739_n9,
         DP_OP_992_186_8739_n8, DP_OP_992_186_8739_n7, DP_OP_987_181_8739_n32,
         DP_OP_987_181_8739_n31, DP_OP_987_181_8739_n30,
         DP_OP_987_181_8739_n29, DP_OP_987_181_8739_n27,
         DP_OP_987_181_8739_n25, DP_OP_987_181_8739_n24,
         DP_OP_987_181_8739_n23, DP_OP_987_181_8739_n21,
         DP_OP_987_181_8739_n20, DP_OP_987_181_8739_n19,
         DP_OP_987_181_8739_n15, DP_OP_987_181_8739_n13,
         DP_OP_987_181_8739_n11, DP_OP_987_181_8739_n9, DP_OP_987_181_8739_n8,
         DP_OP_987_181_8739_n7, DP_OP_981_175_8739_n32, DP_OP_981_175_8739_n31,
         DP_OP_981_175_8739_n30, DP_OP_981_175_8739_n29,
         DP_OP_981_175_8739_n28, DP_OP_981_175_8739_n23,
         DP_OP_981_175_8739_n15, DP_OP_981_175_8739_n13,
         DP_OP_981_175_8739_n11, DP_OP_981_175_8739_n9, DP_OP_981_175_8739_n8,
         DP_OP_981_175_8739_n7, DP_OP_981_175_8739_n5, DP_OP_981_175_8739_n4,
         DP_OP_981_175_8739_n3, DP_OP_981_175_8739_n2, DP_OP_981_175_8739_n1,
         DP_OP_985_179_8739_n31, DP_OP_985_179_8739_n30,
         DP_OP_985_179_8739_n29, DP_OP_985_179_8739_n28,
         DP_OP_985_179_8739_n27, DP_OP_985_179_8739_n25,
         DP_OP_985_179_8739_n24, DP_OP_985_179_8739_n19,
         DP_OP_985_179_8739_n11, DP_OP_985_179_8739_n7, DP_OP_985_179_8739_n3,
         DP_OP_985_179_8739_n2, DP_OP_985_179_8739_n1, DP_OP_983_177_8739_n32,
         DP_OP_983_177_8739_n31, DP_OP_983_177_8739_n30,
         DP_OP_983_177_8739_n29, DP_OP_983_177_8739_n28,
         DP_OP_983_177_8739_n23, DP_OP_983_177_8739_n21,
         DP_OP_983_177_8739_n20, DP_OP_983_177_8739_n19,
         DP_OP_983_177_8739_n17, DP_OP_983_177_8739_n16,
         DP_OP_983_177_8739_n15, DP_OP_983_177_8739_n11, DP_OP_983_177_8739_n9,
         DP_OP_983_177_8739_n8, DP_OP_983_177_8739_n3, DP_OP_983_177_8739_n2,
         DP_OP_983_177_8739_n1, DP_OP_984_178_8739_n28, DP_OP_984_178_8739_n27,
         DP_OP_984_178_8739_n26, DP_OP_984_178_8739_n25,
         DP_OP_984_178_8739_n24, DP_OP_984_178_8739_n23,
         DP_OP_984_178_8739_n19, DP_OP_984_178_8739_n17,
         DP_OP_984_178_8739_n16, DP_OP_984_178_8739_n15,
         DP_OP_984_178_8739_n13, DP_OP_984_178_8739_n12,
         DP_OP_984_178_8739_n11, DP_OP_984_178_8739_n9, DP_OP_984_178_8739_n8,
         DP_OP_984_178_8739_n7, DP_OP_980_174_8739_n28, DP_OP_980_174_8739_n26,
         DP_OP_980_174_8739_n25, DP_OP_980_174_8739_n19,
         DP_OP_980_174_8739_n17, DP_OP_980_174_8739_n16,
         DP_OP_980_174_8739_n15, DP_OP_980_174_8739_n13,
         DP_OP_980_174_8739_n12, DP_OP_980_174_8739_n11, DP_OP_980_174_8739_n9,
         DP_OP_980_174_8739_n8, DP_OP_980_174_8739_n7, DP_OP_988_182_8739_n28,
         DP_OP_988_182_8739_n27, DP_OP_988_182_8739_n26,
         DP_OP_988_182_8739_n25, DP_OP_988_182_8739_n24,
         DP_OP_988_182_8739_n23, DP_OP_988_182_8739_n21,
         DP_OP_988_182_8739_n20, DP_OP_988_182_8739_n19,
         DP_OP_988_182_8739_n17, DP_OP_988_182_8739_n16,
         DP_OP_988_182_8739_n15, DP_OP_988_182_8739_n13,
         DP_OP_988_182_8739_n12, DP_OP_988_182_8739_n11, DP_OP_988_182_8739_n9,
         DP_OP_988_182_8739_n8, DP_OP_988_182_8739_n7, DP_OP_988_182_8739_n3,
         DP_OP_988_182_8739_n2, DP_OP_988_182_8739_n1, DP_OP_982_176_8739_n23,
         DP_OP_982_176_8739_n22, DP_OP_982_176_8739_n21,
         DP_OP_982_176_8739_n19, DP_OP_982_176_8739_n17,
         DP_OP_982_176_8739_n16, DP_OP_982_176_8739_n15,
         DP_OP_982_176_8739_n11, DP_OP_982_176_8739_n9, DP_OP_982_176_8739_n8,
         DP_OP_982_176_8739_n7, DP_OP_986_180_8739_n18, DP_OP_986_180_8739_n17,
         DP_OP_986_180_8739_n15, DP_OP_986_180_8739_n11, DP_OP_986_180_8739_n7,
         DP_OP_982J1_125_6202_n182, DP_OP_982J1_125_6202_n181,
         DP_OP_982J1_125_6202_n180, DP_OP_982J1_125_6202_n177,
         DP_OP_982J1_125_6202_n175, DP_OP_982J1_125_6202_n139,
         DP_OP_982J1_125_6202_n137, DP_OP_982J1_125_6202_n136,
         DP_OP_982J1_125_6202_n135, DP_OP_982J1_125_6202_n132,
         DP_OP_982J1_125_6202_n131, DP_OP_982J1_125_6202_n130,
         DP_OP_982J1_125_6202_n129, DP_OP_982J1_125_6202_n128,
         DP_OP_982J1_125_6202_n127, DP_OP_982J1_125_6202_n124,
         DP_OP_982J1_125_6202_n123, DP_OP_982J1_125_6202_n122,
         DP_OP_982J1_125_6202_n121, DP_OP_982J1_125_6202_n120,
         DP_OP_982J1_125_6202_n119, DP_OP_982J1_125_6202_n117,
         DP_OP_982J1_125_6202_n113, DP_OP_982J1_125_6202_n112,
         DP_OP_982J1_125_6202_n108, DP_OP_982J1_125_6202_n107,
         DP_OP_982J1_125_6202_n105, DP_OP_982J1_125_6202_n104,
         DP_OP_982J1_125_6202_n100, DP_OP_982J1_125_6202_n99,
         DP_OP_982J1_125_6202_n98, DP_OP_982J1_125_6202_n97,
         DP_OP_982J1_125_6202_n96, DP_OP_982J1_125_6202_n95,
         DP_OP_982J1_125_6202_n90, DP_OP_982J1_125_6202_n89,
         DP_OP_982J1_125_6202_n84, DP_OP_982J1_125_6202_n83,
         DP_OP_982J1_125_6202_n78, DP_OP_982J1_125_6202_n77,
         DP_OP_982J1_125_6202_n75, DP_OP_982J1_125_6202_n74,
         DP_OP_982J1_125_6202_n73, DP_OP_982J1_125_6202_n68,
         DP_OP_982J1_125_6202_n67, DP_OP_982J1_125_6202_n66,
         DP_OP_982J1_125_6202_n63, DP_OP_982J1_125_6202_n62,
         DP_OP_982J1_125_6202_n61, DP_OP_982J1_125_6202_n58,
         DP_OP_982J1_125_6202_n57, DP_OP_982J1_125_6202_n56,
         DP_OP_982J1_125_6202_n45, DP_OP_982J1_125_6202_n44,
         DP_OP_982J1_125_6202_n38, DP_OP_982J1_125_6202_n37,
         DP_OP_982J1_125_6202_n35, DP_OP_982J1_125_6202_n34,
         DP_OP_982J1_125_6202_n33, DP_OP_982J1_125_6202_n31,
         DP_OP_982J1_125_6202_n28, DP_OP_982J1_125_6202_n27,
         DP_OP_982J1_125_6202_n24, DP_OP_982J1_125_6202_n20,
         DP_OP_982J1_125_6202_n16, DP_OP_982J1_125_6202_n15,
         DP_OP_982J1_125_6202_n12, DP_OP_982J1_125_6202_n10,
         DP_OP_982J1_125_6202_n9, DP_OP_982J1_125_6202_n8,
         DP_OP_982J1_125_6202_n4, DP_OP_981J1_124_6202_n140,
         DP_OP_981J1_124_6202_n137, DP_OP_981J1_124_6202_n135,
         DP_OP_981J1_124_6202_n131, DP_OP_981J1_124_6202_n129,
         DP_OP_981J1_124_6202_n127, DP_OP_981J1_124_6202_n124,
         DP_OP_981J1_124_6202_n123, DP_OP_981J1_124_6202_n122,
         DP_OP_981J1_124_6202_n121, DP_OP_981J1_124_6202_n120,
         DP_OP_981J1_124_6202_n119, DP_OP_981J1_124_6202_n117,
         DP_OP_981J1_124_6202_n114, DP_OP_981J1_124_6202_n113,
         DP_OP_981J1_124_6202_n112, DP_OP_981J1_124_6202_n109,
         DP_OP_981J1_124_6202_n108, DP_OP_981J1_124_6202_n107,
         DP_OP_981J1_124_6202_n106, DP_OP_981J1_124_6202_n105,
         DP_OP_981J1_124_6202_n104, DP_OP_981J1_124_6202_n101,
         DP_OP_981J1_124_6202_n100, DP_OP_981J1_124_6202_n99,
         DP_OP_981J1_124_6202_n98, DP_OP_981J1_124_6202_n97,
         DP_OP_981J1_124_6202_n96, DP_OP_981J1_124_6202_n95,
         DP_OP_981J1_124_6202_n90, DP_OP_981J1_124_6202_n89,
         DP_OP_981J1_124_6202_n84, DP_OP_981J1_124_6202_n83,
         DP_OP_981J1_124_6202_n78, DP_OP_981J1_124_6202_n77,
         DP_OP_981J1_124_6202_n73, DP_OP_981J1_124_6202_n62,
         DP_OP_981J1_124_6202_n61, DP_OP_981J1_124_6202_n57,
         DP_OP_981J1_124_6202_n45, DP_OP_981J1_124_6202_n44,
         DP_OP_981J1_124_6202_n38, DP_OP_981J1_124_6202_n37,
         DP_OP_981J1_124_6202_n33, DP_OP_981J1_124_6202_n31,
         DP_OP_981J1_124_6202_n24, DP_OP_981J1_124_6202_n20,
         DP_OP_981J1_124_6202_n17, DP_OP_981J1_124_6202_n16,
         DP_OP_981J1_124_6202_n15, DP_OP_981J1_124_6202_n11,
         DP_OP_981J1_124_6202_n10, DP_OP_981J1_124_6202_n9,
         DP_OP_981J1_124_6202_n8, DP_OP_981J1_124_6202_n4, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n104, n106,
         n107, n108, n114, n115, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n209,
         n210, n220, n221, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n275, n276,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n665, n666, n667, n668, n669, n670, n671, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n916, n917, n918,
         n919, n920, n921, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1102, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1469, n1470, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628;
  wire   [2:0] StateMC;
  wire   [3:0] Debug_reg;
  wire   [7:0] Final_Exponent_reg;
  wire   [10:1] Final_Mantissa_reg;

  DFFRX1 Add_sign_reg_reg ( .D(n1103), .CLK(CLK), .CLRB(n73), .Q(n307), .QB(
        n277) );
  DFFRX1 Final_Mantissa_reg_reg_10_ ( .D(n1062), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[10]), .QB(n296) );
  DFFRX1 Final_Exponent_reg_reg_7_ ( .D(n346), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[7]), .QB(n405) );
  DFFRX1 StateMC_reg_1_ ( .D(n922), .CLK(CLK), .CLRB(n73), .Q(n300), .QB(
        StateMC[1]) );
  DFFRX1 Op2_Sign_reg_reg ( .D(n1090), .CLK(CLK), .CLRB(n73), .Q(Op2_Sign_reg), 
        .QB(n306) );
  DFFRX1 G_reg_reg ( .D(n1072), .CLK(CLK), .CLRB(n73), .Q(n189), .QB(
        add_x_35_A_2_) );
  DFFRX1 Final_Mantissa_reg_reg_2_ ( .D(n664), .CLK(CLK), .CLRB(n73), .Q(n312), 
        .QB(Final_Mantissa_reg[2]) );
  DFFRX1 Final_Mantissa_reg_reg_1_ ( .D(n672), .CLK(CLK), .CLRB(n73), .Q(n299), 
        .QB(Final_Mantissa_reg[1]) );
  DFFRX1 Final_Mantissa_reg_reg_0_ ( .D(n113), .CLK(CLK), .CLRB(n73), .Q(N691), 
        .QB(n297) );
  DFFRX1 Final_Mantissa_reg_reg_8_ ( .D(n1064), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[8]), .QB(n314) );
  DFFRX1 exc_reg_reg_0_ ( .D(n1092), .CLK(CLK), .CLRB(n73), .Q(exc_reg_0_), 
        .QB(n317) );
  DFFRX1 StateMC_reg_0_ ( .D(n991), .CLK(CLK), .CLRB(n73), .Q(n301), .QB(
        StateMC[0]) );
  DFFRX1 StateMC_reg_2_ ( .D(n915), .CLK(CLK), .CLRB(n73), .Q(n313), .QB(
        StateMC[2]) );
  DFFRX1 Op1_Sign_reg_reg ( .D(n1081), .CLK(CLK), .CLRB(n73), .Q(Op1_Sign_reg), 
        .QB(n305) );
  DFFRX1 Op1_Mantissa_reg_reg_6_ ( .D(n1083), .CLK(CLK), .CLRB(n73), .QB(n213)
         );
  DFFRX1 Op1_Mantissa_reg_reg_5_ ( .D(n1084), .CLK(CLK), .CLRB(n73), .QB(n214)
         );
  DFFRX1 Op1_Mantissa_reg_reg_4_ ( .D(n1085), .CLK(CLK), .CLRB(n73), .QB(n215)
         );
  DFFRX1 Op1_Mantissa_reg_reg_3_ ( .D(n1086), .CLK(CLK), .CLRB(n73), .QB(n216)
         );
  DFFRX1 Op1_Mantissa_reg_reg_2_ ( .D(n1087), .CLK(CLK), .CLRB(n73), .QB(n217)
         );
  DFFRX1 Op1_Mantissa_reg_reg_1_ ( .D(n1088), .CLK(CLK), .CLRB(n73), .QB(n218)
         );
  DFFRX1 Op1_Mantissa_reg_reg_0_ ( .D(n1089), .CLK(CLK), .CLRB(n73), .QB(n219)
         );
  DFFRX1 Op2_Mantissa_reg_reg_7_ ( .D(n1073), .CLK(CLK), .CLRB(n73), .Q(
        Op2_Mantissa_reg_7_), .QB(n321) );
  DFFRX1 R_reg_reg ( .D(n1070), .CLK(CLK), .CLRB(n73), .Q(n861), .QB(
        add_x_35_A_1_) );
  DFFRX1 S_reg_reg ( .D(n1071), .CLK(CLK), .CLRB(n73), .Q(n188), .QB(
        add_x_35_A_0_) );
  DFFRX1 Adder_datain2_reg_8_ ( .D(n124), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[8]) );
  DFFRX1 Adder_datain2_reg_7_ ( .D(n123), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[7]) );
  DFFRX1 Adder_datain1_reg_6_ ( .D(N258), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[6]) );
  DFFRX1 Adder_datain1_reg_5_ ( .D(N257), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[5]) );
  DFFRX1 Adder_datain1_reg_4_ ( .D(N256), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[4]) );
  DFFRX1 Adder_datain1_reg_3_ ( .D(N255), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[3]) );
  DFFRX1 Adder_datain1_reg_2_ ( .D(N254), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[2]) );
  DFFRX1 Adder_datain1_reg_1_ ( .D(N253), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[1]) );
  DFFRX1 Adder_datain1_reg_0_ ( .D(N252), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[0]) );
  DFFRX1 carry_reg_reg ( .D(n1061), .CLK(CLK), .CLRB(n73), .Q(carry_reg), .QB(
        n303) );
  DFFRX1 Final_Mantissa_reg_reg_9_ ( .D(n1063), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[9]), .QB(n310) );
  DFFRX1 Final_Mantissa_reg_reg_7_ ( .D(n1065), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[7]), .QB(n309) );
  DFFRX1 Final_Mantissa_reg_reg_6_ ( .D(n1066), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[6]), .QB(n186) );
  DFFRX1 Final_Mantissa_reg_reg_5_ ( .D(n1067), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[5]), .QB(n311) );
  DFFRX1 Final_Mantissa_reg_reg_4_ ( .D(n1068), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[4]), .QB(n298) );
  DFFRX1 Final_Mantissa_reg_reg_3_ ( .D(n1069), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[3]), .QB(n308) );
  DFFRX1 Debug_valid_reg_reg ( .D(n103), .CLK(CLK), .CLRB(n73), .Q(
        Debug_valid_reg), .QB(n323) );
  DFFRX1 Adder_valid_reg ( .D(n1091), .CLK(CLK), .CLRB(n73), .Q(Adder_valid), 
        .QB(n322) );
  DFFRX1 exc_reg_reg_1_ ( .D(n1093), .CLK(CLK), .CLRB(n73), .Q(n320), .QB(n223) );
  DFFRX1 exc_reg_reg_2_ ( .D(n1101), .CLK(CLK), .CLRB(n73), .Q(n302), .QB(n222) );
  DFFRX1 Final_Sign_reg_reg ( .D(n1060), .CLK(CLK), .CLRB(n73), .Q(n324), .QB(
        n274) );
  DFFRX1 Op1_Mantissa_reg_reg_7_ ( .D(n1082), .CLK(CLK), .CLRB(n73), .QB(n212)
         );
  DFFRX1 Adder_datain1_reg_7_ ( .D(N259), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[7]) );
  DFFRX1 Op2_Mantissa_reg_reg_0_ ( .D(n1080), .CLK(CLK), .CLRB(n73), .Q(n1477), 
        .QB(add_x_35_A_3_) );
  DFFRX1 Adder_datain2_reg_0_ ( .D(n116), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[0]) );
  DFFRX1 Op2_Mantissa_reg_reg_1_ ( .D(n1079), .CLK(CLK), .CLRB(n73), .Q(n1552), 
        .QB(add_x_35_A_4_) );
  DFFRX1 Adder_datain2_reg_1_ ( .D(n117), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[1]) );
  DFFRX1 Op2_Mantissa_reg_reg_2_ ( .D(n1078), .CLK(CLK), .CLRB(n73), .Q(n1554), 
        .QB(add_x_35_A_5_) );
  DFFRX1 Adder_datain2_reg_2_ ( .D(n118), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[2]) );
  DFFRX1 Op2_Mantissa_reg_reg_3_ ( .D(n1077), .CLK(CLK), .CLRB(n73), .Q(n315), 
        .QB(add_x_35_A_6_) );
  DFFRX1 Adder_datain2_reg_3_ ( .D(n119), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[3]) );
  DFFRX1 Op2_Mantissa_reg_reg_4_ ( .D(n1076), .CLK(CLK), .CLRB(n73), .Q(n316), 
        .QB(add_x_35_A_7_) );
  DFFRX1 Adder_datain2_reg_4_ ( .D(n120), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[4]) );
  DFFRX1 Op2_Mantissa_reg_reg_5_ ( .D(n1075), .CLK(CLK), .CLRB(n73), .Q(n318), 
        .QB(add_x_35_A_8_) );
  DFFRX1 Adder_datain2_reg_5_ ( .D(n121), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[5]) );
  DFFRX1 Op2_Mantissa_reg_reg_6_ ( .D(n1074), .CLK(CLK), .CLRB(n73), .Q(n319), 
        .QB(add_x_35_A_9_) );
  DFFRX1 Adder_datain2_reg_6_ ( .D(n122), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[6]) );
  DFFRX1 Final_Exponent_reg_reg_0_ ( .D(n1094), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[0]), .QB(n292) );
  DFFRX1 Final_Exponent_reg_reg_1_ ( .D(n1095), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[1]), .QB(n406) );
  DFFRX1 Final_Exponent_reg_reg_2_ ( .D(n1096), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[2]), .QB(n293) );
  DFFRX1 Final_Exponent_reg_reg_3_ ( .D(n1097), .CLK(CLK), .CLRB(n73), .Q(n185), .QB(n294) );
  DFFRX1 Final_Exponent_reg_reg_4_ ( .D(n1098), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[4]), .QB(n408) );
  DFFRX1 Final_Exponent_reg_reg_5_ ( .D(n1099), .CLK(CLK), .CLRB(n73), .Q(n187), .QB(n304) );
  DFFRX1 Final_Exponent_reg_reg_6_ ( .D(n1100), .CLK(CLK), .CLRB(n73), .QB(
        n295) );
  DFFRX1 ExcCheck_valid_reg ( .D(N270), .CLK(CLK), .CLRB(n73), .Q(
        ExcCheck_valid) );
  DFFRX1 Debug_reg_reg_3_ ( .D(n112), .CLK(CLK), .CLRB(n73), .Q(Debug_reg[3])
         );
  DFFRX1 Debug_reg_reg_2_ ( .D(n111), .CLK(CLK), .CLRB(n73), .Q(Debug_reg[2])
         );
  DFFRX1 Debug_reg_reg_1_ ( .D(n110), .CLK(CLK), .CLRB(n73), .Q(Debug_reg[1])
         );
  DFFRX1 Debug_reg_reg_0_ ( .D(n109), .CLK(CLK), .CLRB(n73), .Q(Debug_reg[0])
         );
  NOR2X1 DP_OP_979_173_2805_U57 ( .IN1(n407), .IN2(n398), .OUT(
        DP_OP_979_173_2805_n55) );
  NOR2X1 DP_OP_979_173_2805_U49 ( .IN1(n407), .IN2(n411), .OUT(
        DP_OP_979_173_2805_n52) );
  NAND2X1 DP_OP_979_173_2805_U47 ( .IN1(DP_OP_979_173_2805_n55), .IN2(n411), 
        .OUT(DP_OP_979_173_2805_n20) );
  NAND2X1 DP_OP_979_173_2805_U45 ( .IN1(n411), .IN2(DP_OP_979_173_2805_n20), 
        .OUT(DP_OP_979_173_2805_n18) );
  NOR2X1 DP_OP_979_173_2805_U40 ( .IN1(DP_OP_979_173_2805_n76), .IN2(
        DP_OP_979_173_2805_n1), .OUT(DP_OP_979_173_2805_n48) );
  NOR2X1 DP_OP_979_173_2805_U39 ( .IN1(DP_OP_979_173_2805_n1), .IN2(n185), 
        .OUT(DP_OP_979_173_2805_n17) );
  NOR2X1 DP_OP_979_173_2805_U38 ( .IN1(DP_OP_979_173_2805_n1), .IN2(
        DP_OP_979_173_2805_n17), .OUT(DP_OP_979_173_2805_n16) );
  NOR2X1 DP_OP_979_173_2805_U37 ( .IN1(DP_OP_979_173_2805_n76), .IN2(
        DP_OP_979_173_2805_n17), .OUT(DP_OP_979_173_2805_n15) );
  NOR2X1 DP_OP_979_173_2805_U36 ( .IN1(DP_OP_979_173_2805_n16), .IN2(
        DP_OP_979_173_2805_n15), .OUT(C1_DATA1_3) );
  NOR2X1 DP_OP_979_173_2805_U32 ( .IN1(DP_OP_979_173_2805_n76), .IN2(
        DP_OP_979_173_2805_n77), .OUT(DP_OP_979_173_2805_n45) );
  NOR2X1 DP_OP_979_173_2805_U30 ( .IN1(DP_OP_979_173_2805_n44), .IN2(
        DP_OP_979_173_2805_n1), .OUT(DP_OP_979_173_2805_n43) );
  NAND2X1 DP_OP_979_173_2805_U28 ( .IN1(DP_OP_979_173_2805_n48), .IN2(
        DP_OP_979_173_2805_n14), .OUT(DP_OP_979_173_2805_n13) );
  NAND2X1 DP_OP_979_173_2805_U21 ( .IN1(DP_OP_979_173_2805_n45), .IN2(n199), 
        .OUT(DP_OP_979_173_2805_n39) );
  NAND2X1 DP_OP_979_173_2805_U18 ( .IN1(DP_OP_979_173_2805_n43), .IN2(
        DP_OP_979_173_2805_n11), .OUT(DP_OP_979_173_2805_n10) );
  NOR2X1 DP_OP_979_173_2805_U12 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_979_173_2805_n79), .OUT(DP_OP_979_173_2805_n35) );
  NOR2X1 DP_OP_989_183_2805_U64 ( .IN1(n919), .IN2(n201), .OUT(
        DP_OP_989_183_2805_n26) );
  NOR2X1 DP_OP_989_183_2805_U63 ( .IN1(n410), .IN2(n201), .OUT(
        DP_OP_989_183_2805_n25) );
  NOR2X1 DP_OP_989_183_2805_U62 ( .IN1(DP_OP_989_183_2805_n26), .IN2(
        DP_OP_989_183_2805_n25), .OUT(C1_DATA11_0) );
  NOR2X1 DP_OP_989_183_2805_U57 ( .IN1(n407), .IN2(n395), .OUT(
        DP_OP_989_183_2805_n55) );
  NOR2X1 DP_OP_989_183_2805_U40 ( .IN1(n185), .IN2(DP_OP_989_183_2805_n1), 
        .OUT(DP_OP_989_183_2805_n48) );
  NOR2X1 DP_OP_989_183_2805_U30 ( .IN1(DP_OP_979_173_2805_n44), .IN2(
        DP_OP_989_183_2805_n1), .OUT(DP_OP_989_183_2805_n43) );
  NOR2X1 DP_OP_989_183_2805_U20 ( .IN1(DP_OP_989_183_2805_n1), .IN2(
        DP_OP_979_173_2805_n39), .OUT(DP_OP_989_183_2805_n38) );
  NAND2X1 DP_OP_989_183_2805_U18 ( .IN1(DP_OP_989_183_2805_n43), .IN2(
        DP_OP_989_183_2805_n11), .OUT(DP_OP_989_183_2805_n10) );
  NOR2X1 DP_OP_989_183_2805_U10 ( .IN1(DP_OP_989_183_2805_n1), .IN2(
        DP_OP_990_184_2805_n34), .OUT(DP_OP_989_183_2805_n2) );
  NAND2X1 DP_OP_989_183_2805_U4 ( .IN1(DP_OP_989_183_2805_n2), .IN2(
        DP_OP_989_183_2805_n5), .OUT(DP_OP_989_183_2805_n4) );
  NOR2X1 DP_OP_990_184_2805_U66 ( .IN1(n410), .IN2(n919), .OUT(
        DP_OP_990_184_2805_n58) );
  NOR2X1 DP_OP_990_184_2805_U64 ( .IN1(n919), .IN2(DP_OP_990_184_2805_n58), 
        .OUT(DP_OP_990_184_2805_n26) );
  NOR2X1 DP_OP_990_184_2805_U63 ( .IN1(n410), .IN2(DP_OP_990_184_2805_n58), 
        .OUT(DP_OP_990_184_2805_n25) );
  NOR2X1 DP_OP_990_184_2805_U62 ( .IN1(DP_OP_990_184_2805_n26), .IN2(
        DP_OP_990_184_2805_n25), .OUT(C1_DATA12_0) );
  NAND2X1 DP_OP_990_184_2805_U56 ( .IN1(DP_OP_990_184_2805_n58), .IN2(n407), 
        .OUT(DP_OP_990_184_2805_n23) );
  NAND2X1 DP_OP_990_184_2805_U55 ( .IN1(DP_OP_990_184_2805_n58), .IN2(
        DP_OP_990_184_2805_n23), .OUT(DP_OP_990_184_2805_n22) );
  NOR2X1 DP_OP_990_184_2805_U40 ( .IN1(DP_OP_979_173_2805_n76), .IN2(
        DP_OP_990_184_2805_n51), .OUT(DP_OP_990_184_2805_n48) );
  NOR2X1 DP_OP_990_184_2805_U30 ( .IN1(DP_OP_979_173_2805_n44), .IN2(
        DP_OP_990_184_2805_n51), .OUT(DP_OP_990_184_2805_n43) );
  NAND2X1 DP_OP_990_184_2805_U28 ( .IN1(DP_OP_990_184_2805_n48), .IN2(
        DP_OP_990_184_2805_n14), .OUT(DP_OP_990_184_2805_n13) );
  NAND2X1 DP_OP_990_184_2805_U19 ( .IN1(DP_OP_990_184_2805_n43), .IN2(n187), 
        .OUT(DP_OP_990_184_2805_n11) );
  NAND2X1 DP_OP_990_184_2805_U18 ( .IN1(DP_OP_990_184_2805_n43), .IN2(
        DP_OP_990_184_2805_n11), .OUT(DP_OP_990_184_2805_n10) );
  NOR2X1 DP_OP_990_184_2805_U10 ( .IN1(DP_OP_990_184_2805_n51), .IN2(
        DP_OP_990_184_2805_n34), .OUT(DP_OP_990_184_2805_n2) );
  NOR2X1 DP_OP_991_185_2805_U62 ( .IN1(DP_OP_989_183_2805_n26), .IN2(
        DP_OP_989_183_2805_n25), .OUT(C1_DATA13_0) );
  NOR2X1 DP_OP_991_185_2805_U40 ( .IN1(n185), .IN2(DP_OP_989_183_2805_n1), 
        .OUT(DP_OP_991_185_2805_n48) );
  NOR2X1 DP_OP_991_185_2805_U30 ( .IN1(DP_OP_979_173_2805_n44), .IN2(
        DP_OP_989_183_2805_n1), .OUT(DP_OP_991_185_2805_n43) );
  NOR2X1 DP_OP_991_185_2805_U20 ( .IN1(DP_OP_989_183_2805_n1), .IN2(
        DP_OP_979_173_2805_n39), .OUT(DP_OP_991_185_2805_n38) );
  NAND2X1 DP_OP_991_185_2805_U18 ( .IN1(DP_OP_991_185_2805_n43), .IN2(
        DP_OP_991_185_2805_n11), .OUT(DP_OP_991_185_2805_n10) );
  NOR2X1 DP_OP_991_185_2805_U10 ( .IN1(DP_OP_989_183_2805_n1), .IN2(
        DP_OP_990_184_2805_n34), .OUT(DP_OP_991_185_2805_n2) );
  NAND2X1 DP_OP_991_185_2805_U4 ( .IN1(DP_OP_991_185_2805_n2), .IN2(
        DP_OP_991_185_2805_n5), .OUT(DP_OP_991_185_2805_n4) );
  NOR2X1 DP_OP_987_181_8739_U40 ( .IN1(Final_Exponent_reg[1]), .IN2(
        Final_Exponent_reg[0]), .OUT(DP_OP_987_181_8739_n27) );
  NOR2X1 DP_OP_987_181_8739_U37 ( .IN1(n410), .IN2(DP_OP_987_181_8739_n27), 
        .OUT(DP_OP_987_181_8739_n25) );
  NOR2X1 DP_OP_987_181_8739_U36 ( .IN1(n407), .IN2(DP_OP_987_181_8739_n27), 
        .OUT(DP_OP_987_181_8739_n24) );
  NOR2X1 DP_OP_987_181_8739_U35 ( .IN1(DP_OP_987_181_8739_n25), .IN2(
        DP_OP_987_181_8739_n24), .OUT(C1_DATA9_1) );
  NOR2X1 DP_OP_987_181_8739_U34 ( .IN1(n411), .IN2(n205), .OUT(
        DP_OP_987_181_8739_n23) );
  NOR2X1 DP_OP_987_181_8739_U31 ( .IN1(n205), .IN2(DP_OP_987_181_8739_n23), 
        .OUT(DP_OP_987_181_8739_n21) );
  NOR2X1 DP_OP_987_181_8739_U30 ( .IN1(n411), .IN2(DP_OP_987_181_8739_n23), 
        .OUT(DP_OP_987_181_8739_n20) );
  NOR2X1 DP_OP_987_181_8739_U29 ( .IN1(DP_OP_987_181_8739_n21), .IN2(
        DP_OP_987_181_8739_n20), .OUT(C1_DATA9_2) );
  NOR2X1 DP_OP_987_181_8739_U19 ( .IN1(DP_OP_987_181_8739_n31), .IN2(
        DP_OP_987_181_8739_n15), .OUT(DP_OP_987_181_8739_n13) );
  NOR2X1 DP_OP_987_181_8739_U13 ( .IN1(DP_OP_987_181_8739_n30), .IN2(
        DP_OP_987_181_8739_n11), .OUT(DP_OP_987_181_8739_n9) );
  NOR2X1 DP_OP_987_181_8739_U12 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_987_181_8739_n11), .OUT(DP_OP_987_181_8739_n8) );
  NOR2X1 DP_OP_987_181_8739_U11 ( .IN1(DP_OP_987_181_8739_n9), .IN2(
        DP_OP_987_181_8739_n8), .OUT(C1_DATA9_5) );
  NOR2X1 DP_OP_987_181_8739_U10 ( .IN1(DP_OP_979_173_2805_n79), .IN2(
        DP_OP_987_181_8739_n29), .OUT(DP_OP_987_181_8739_n7) );
  NOR2X1 DP_OP_981_175_8739_U19 ( .IN1(DP_OP_981_175_8739_n31), .IN2(
        DP_OP_981_175_8739_n15), .OUT(DP_OP_981_175_8739_n13) );
  NOR2X1 DP_OP_981_175_8739_U13 ( .IN1(DP_OP_981_175_8739_n30), .IN2(
        DP_OP_981_175_8739_n11), .OUT(DP_OP_981_175_8739_n9) );
  NOR2X1 DP_OP_981_175_8739_U12 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_981_175_8739_n11), .OUT(DP_OP_981_175_8739_n8) );
  NOR2X1 DP_OP_981_175_8739_U11 ( .IN1(DP_OP_981_175_8739_n9), .IN2(
        DP_OP_981_175_8739_n8), .OUT(C1_DATA3_5) );
  NOR2X1 DP_OP_981_175_8739_U10 ( .IN1(DP_OP_979_173_2805_n79), .IN2(
        DP_OP_981_175_8739_n29), .OUT(DP_OP_981_175_8739_n7) );
  NOR2X1 DP_OP_981_175_8739_U7 ( .IN1(DP_OP_981_175_8739_n29), .IN2(
        DP_OP_981_175_8739_n7), .OUT(DP_OP_981_175_8739_n5) );
  NOR2X1 DP_OP_981_175_8739_U6 ( .IN1(DP_OP_979_173_2805_n79), .IN2(
        DP_OP_981_175_8739_n7), .OUT(DP_OP_981_175_8739_n4) );
  NOR2X1 DP_OP_981_175_8739_U5 ( .IN1(DP_OP_981_175_8739_n5), .IN2(
        DP_OP_981_175_8739_n4), .OUT(C1_DATA3_6) );
  NOR2X1 DP_OP_981_175_8739_U4 ( .IN1(DP_OP_981_175_8739_n28), .IN2(
        DP_OP_979_173_2805_n80), .OUT(DP_OP_981_175_8739_n3) );
  NOR2X1 DP_OP_981_175_8739_U3 ( .IN1(DP_OP_981_175_8739_n28), .IN2(
        DP_OP_981_175_8739_n3), .OUT(DP_OP_981_175_8739_n2) );
  NOR2X1 DP_OP_981_175_8739_U2 ( .IN1(DP_OP_979_173_2805_n80), .IN2(
        DP_OP_981_175_8739_n3), .OUT(DP_OP_981_175_8739_n1) );
  NOR2X1 DP_OP_981_175_8739_U1 ( .IN1(DP_OP_981_175_8739_n2), .IN2(
        DP_OP_981_175_8739_n1), .OUT(C1_DATA3_7) );
  NOR2X1 DP_OP_985_179_8739_U16 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_985_179_8739_n30), .OUT(DP_OP_985_179_8739_n11) );
  NOR2X1 DP_OP_985_179_8739_U10 ( .IN1(DP_OP_979_173_2805_n79), .IN2(
        DP_OP_985_179_8739_n29), .OUT(DP_OP_985_179_8739_n7) );
  NOR2X1 DP_OP_985_179_8739_U4 ( .IN1(DP_OP_985_179_8739_n28), .IN2(
        DP_OP_979_173_2805_n80), .OUT(DP_OP_985_179_8739_n3) );
  NOR2X1 DP_OP_985_179_8739_U3 ( .IN1(DP_OP_985_179_8739_n28), .IN2(
        DP_OP_985_179_8739_n3), .OUT(DP_OP_985_179_8739_n2) );
  NOR2X1 DP_OP_985_179_8739_U2 ( .IN1(DP_OP_979_173_2805_n80), .IN2(
        DP_OP_985_179_8739_n3), .OUT(DP_OP_985_179_8739_n1) );
  NOR2X1 DP_OP_985_179_8739_U1 ( .IN1(DP_OP_985_179_8739_n2), .IN2(
        DP_OP_985_179_8739_n1), .OUT(C1_DATA7_7) );
  NOR2X1 DP_OP_983_177_8739_U35 ( .IN1(DP_OP_987_181_8739_n25), .IN2(
        DP_OP_987_181_8739_n24), .OUT(C1_DATA5_1) );
  NOR2X1 DP_OP_983_177_8739_U28 ( .IN1(n185), .IN2(DP_OP_983_177_8739_n32), 
        .OUT(DP_OP_983_177_8739_n19) );
  NOR2X1 DP_OP_983_177_8739_U25 ( .IN1(DP_OP_983_177_8739_n32), .IN2(
        DP_OP_983_177_8739_n19), .OUT(DP_OP_983_177_8739_n17) );
  NOR2X1 DP_OP_983_177_8739_U24 ( .IN1(DP_OP_979_173_2805_n76), .IN2(
        DP_OP_983_177_8739_n19), .OUT(DP_OP_983_177_8739_n16) );
  NOR2X1 DP_OP_983_177_8739_U23 ( .IN1(DP_OP_983_177_8739_n17), .IN2(
        DP_OP_983_177_8739_n16), .OUT(C1_DATA5_3) );
  NOR2X1 DP_OP_983_177_8739_U22 ( .IN1(DP_OP_979_173_2805_n77), .IN2(
        DP_OP_983_177_8739_n31), .OUT(DP_OP_983_177_8739_n15) );
  NOR2X1 DP_OP_983_177_8739_U13 ( .IN1(DP_OP_983_177_8739_n30), .IN2(
        DP_OP_983_177_8739_n11), .OUT(DP_OP_983_177_8739_n9) );
  NOR2X1 DP_OP_983_177_8739_U12 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_983_177_8739_n11), .OUT(DP_OP_983_177_8739_n8) );
  NOR2X1 DP_OP_983_177_8739_U11 ( .IN1(DP_OP_983_177_8739_n9), .IN2(
        DP_OP_983_177_8739_n8), .OUT(C1_DATA5_5) );
  NOR2X1 DP_OP_983_177_8739_U4 ( .IN1(DP_OP_983_177_8739_n28), .IN2(
        DP_OP_979_173_2805_n80), .OUT(DP_OP_983_177_8739_n3) );
  NOR2X1 DP_OP_983_177_8739_U3 ( .IN1(DP_OP_983_177_8739_n28), .IN2(
        DP_OP_983_177_8739_n3), .OUT(DP_OP_983_177_8739_n2) );
  NOR2X1 DP_OP_983_177_8739_U2 ( .IN1(DP_OP_979_173_2805_n80), .IN2(
        DP_OP_983_177_8739_n3), .OUT(DP_OP_983_177_8739_n1) );
  NOR2X1 DP_OP_983_177_8739_U1 ( .IN1(DP_OP_983_177_8739_n2), .IN2(
        DP_OP_983_177_8739_n1), .OUT(C1_DATA5_7) );
  NOR2X1 DP_OP_984_178_8739_U25 ( .IN1(DP_OP_984_178_8739_n28), .IN2(
        DP_OP_984_178_8739_n19), .OUT(DP_OP_984_178_8739_n17) );
  NOR2X1 DP_OP_984_178_8739_U24 ( .IN1(n185), .IN2(DP_OP_984_178_8739_n19), 
        .OUT(DP_OP_984_178_8739_n16) );
  NOR2X1 DP_OP_984_178_8739_U23 ( .IN1(DP_OP_984_178_8739_n17), .IN2(
        DP_OP_984_178_8739_n16), .OUT(C1_DATA6_3) );
  NOR2X1 DP_OP_984_178_8739_U19 ( .IN1(DP_OP_984_178_8739_n27), .IN2(
        DP_OP_984_178_8739_n15), .OUT(DP_OP_984_178_8739_n13) );
  NOR2X1 DP_OP_984_178_8739_U18 ( .IN1(DP_OP_979_173_2805_n77), .IN2(
        DP_OP_984_178_8739_n15), .OUT(DP_OP_984_178_8739_n12) );
  NOR2X1 DP_OP_984_178_8739_U17 ( .IN1(DP_OP_984_178_8739_n13), .IN2(
        DP_OP_984_178_8739_n12), .OUT(C1_DATA6_4) );
  NOR2X1 DP_OP_984_178_8739_U16 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_984_178_8739_n26), .OUT(DP_OP_984_178_8739_n11) );
  NOR2X1 DP_OP_984_178_8739_U13 ( .IN1(DP_OP_984_178_8739_n26), .IN2(
        DP_OP_984_178_8739_n11), .OUT(DP_OP_984_178_8739_n9) );
  NOR2X1 DP_OP_984_178_8739_U12 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_984_178_8739_n11), .OUT(DP_OP_984_178_8739_n8) );
  NOR2X1 DP_OP_984_178_8739_U11 ( .IN1(DP_OP_984_178_8739_n9), .IN2(
        DP_OP_984_178_8739_n8), .OUT(C1_DATA6_5) );
  NOR2X1 DP_OP_984_178_8739_U10 ( .IN1(DP_OP_979_173_2805_n79), .IN2(
        DP_OP_984_178_8739_n25), .OUT(DP_OP_984_178_8739_n7) );
  NOR2X1 DP_OP_980_174_8739_U25 ( .IN1(DP_OP_980_174_8739_n28), .IN2(
        DP_OP_980_174_8739_n19), .OUT(DP_OP_980_174_8739_n17) );
  NOR2X1 DP_OP_980_174_8739_U24 ( .IN1(DP_OP_979_173_2805_n76), .IN2(
        DP_OP_980_174_8739_n19), .OUT(DP_OP_980_174_8739_n16) );
  NOR2X1 DP_OP_980_174_8739_U23 ( .IN1(DP_OP_980_174_8739_n17), .IN2(
        DP_OP_980_174_8739_n16), .OUT(C1_DATA2_3) );
  NOR2X1 DP_OP_980_174_8739_U22 ( .IN1(DP_OP_979_173_2805_n77), .IN2(n397), 
        .OUT(DP_OP_980_174_8739_n15) );
  NOR2X1 DP_OP_980_174_8739_U19 ( .IN1(n397), .IN2(DP_OP_980_174_8739_n15), 
        .OUT(DP_OP_980_174_8739_n13) );
  NOR2X1 DP_OP_980_174_8739_U18 ( .IN1(DP_OP_979_173_2805_n77), .IN2(
        DP_OP_980_174_8739_n15), .OUT(DP_OP_980_174_8739_n12) );
  NOR2X1 DP_OP_980_174_8739_U17 ( .IN1(DP_OP_980_174_8739_n13), .IN2(
        DP_OP_980_174_8739_n12), .OUT(C1_DATA2_4) );
  NOR2X1 DP_OP_980_174_8739_U16 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_980_174_8739_n26), .OUT(DP_OP_980_174_8739_n11) );
  NOR2X1 DP_OP_980_174_8739_U13 ( .IN1(DP_OP_980_174_8739_n26), .IN2(
        DP_OP_980_174_8739_n11), .OUT(DP_OP_980_174_8739_n9) );
  NOR2X1 DP_OP_980_174_8739_U12 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_980_174_8739_n11), .OUT(DP_OP_980_174_8739_n8) );
  NOR2X1 DP_OP_980_174_8739_U11 ( .IN1(DP_OP_980_174_8739_n9), .IN2(
        DP_OP_980_174_8739_n8), .OUT(C1_DATA2_5) );
  NOR2X1 DP_OP_980_174_8739_U10 ( .IN1(DP_OP_979_173_2805_n79), .IN2(
        DP_OP_980_174_8739_n25), .OUT(DP_OP_980_174_8739_n7) );
  NOR2X1 DP_OP_988_182_8739_U34 ( .IN1(n411), .IN2(n407), .OUT(
        DP_OP_988_182_8739_n23) );
  NOR2X1 DP_OP_988_182_8739_U31 ( .IN1(n407), .IN2(DP_OP_988_182_8739_n23), 
        .OUT(DP_OP_988_182_8739_n21) );
  NOR2X1 DP_OP_988_182_8739_U30 ( .IN1(n411), .IN2(DP_OP_988_182_8739_n23), 
        .OUT(DP_OP_988_182_8739_n20) );
  NOR2X1 DP_OP_988_182_8739_U29 ( .IN1(DP_OP_988_182_8739_n21), .IN2(
        DP_OP_988_182_8739_n20), .OUT(C1_DATA10_2) );
  NOR2X1 DP_OP_988_182_8739_U19 ( .IN1(DP_OP_988_182_8739_n27), .IN2(
        DP_OP_988_182_8739_n15), .OUT(DP_OP_988_182_8739_n13) );
  NOR2X1 DP_OP_988_182_8739_U18 ( .IN1(DP_OP_979_173_2805_n77), .IN2(
        DP_OP_988_182_8739_n15), .OUT(DP_OP_988_182_8739_n12) );
  NOR2X1 DP_OP_988_182_8739_U13 ( .IN1(DP_OP_988_182_8739_n26), .IN2(
        DP_OP_988_182_8739_n11), .OUT(DP_OP_988_182_8739_n9) );
  NOR2X1 DP_OP_988_182_8739_U12 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_988_182_8739_n11), .OUT(DP_OP_988_182_8739_n8) );
  NOR2X1 DP_OP_988_182_8739_U11 ( .IN1(DP_OP_988_182_8739_n9), .IN2(
        DP_OP_988_182_8739_n8), .OUT(C1_DATA10_5) );
  NOR2X1 DP_OP_988_182_8739_U10 ( .IN1(DP_OP_979_173_2805_n79), .IN2(
        DP_OP_988_182_8739_n25), .OUT(DP_OP_988_182_8739_n7) );
  NOR2X1 DP_OP_988_182_8739_U4 ( .IN1(DP_OP_988_182_8739_n24), .IN2(
        DP_OP_979_173_2805_n80), .OUT(DP_OP_988_182_8739_n3) );
  NOR2X1 DP_OP_988_182_8739_U3 ( .IN1(DP_OP_988_182_8739_n24), .IN2(
        DP_OP_988_182_8739_n3), .OUT(DP_OP_988_182_8739_n2) );
  NOR2X1 DP_OP_988_182_8739_U2 ( .IN1(DP_OP_979_173_2805_n80), .IN2(
        DP_OP_988_182_8739_n3), .OUT(DP_OP_988_182_8739_n1) );
  NOR2X1 DP_OP_988_182_8739_U1 ( .IN1(DP_OP_988_182_8739_n2), .IN2(
        DP_OP_988_182_8739_n1), .OUT(C1_DATA10_7) );
  NOR2X1 DP_OP_982_176_8739_U25 ( .IN1(n185), .IN2(DP_OP_982_176_8739_n19), 
        .OUT(DP_OP_982_176_8739_n17) );
  NOR2X1 DP_OP_982_176_8739_U24 ( .IN1(n411), .IN2(DP_OP_982_176_8739_n19), 
        .OUT(DP_OP_982_176_8739_n16) );
  NOR2X1 DP_OP_982_176_8739_U23 ( .IN1(DP_OP_982_176_8739_n17), .IN2(
        DP_OP_982_176_8739_n16), .OUT(C1_DATA4_3) );
  NOR2X1 DP_OP_982_176_8739_U16 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_982_176_8739_n22), .OUT(DP_OP_982_176_8739_n11) );
  NOR2X1 DP_OP_982_176_8739_U13 ( .IN1(DP_OP_982_176_8739_n22), .IN2(
        DP_OP_982_176_8739_n11), .OUT(DP_OP_982_176_8739_n9) );
  NOR2X1 DP_OP_982_176_8739_U12 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_982_176_8739_n11), .OUT(DP_OP_982_176_8739_n8) );
  NOR2X1 DP_OP_982_176_8739_U11 ( .IN1(DP_OP_982_176_8739_n9), .IN2(
        DP_OP_982_176_8739_n8), .OUT(C1_DATA4_5) );
  NOR2X1 DP_OP_982_176_8739_U10 ( .IN1(DP_OP_979_173_2805_n79), .IN2(
        DP_OP_982_176_8739_n21), .OUT(DP_OP_982_176_8739_n7) );
  NOR2X1 DP_OP_986_180_8739_U22 ( .IN1(DP_OP_979_173_2805_n77), .IN2(n185), 
        .OUT(DP_OP_986_180_8739_n15) );
  NOR2X1 DP_OP_986_180_8739_U16 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_986_180_8739_n18), .OUT(DP_OP_986_180_8739_n11) );
  NOR2X1 DP_OP_986_180_8739_U10 ( .IN1(DP_OP_979_173_2805_n79), .IN2(
        DP_OP_986_180_8739_n17), .OUT(DP_OP_986_180_8739_n7) );
  NAND2X1 DP_OP_992_186_8739_U24 ( .IN1(DP_OP_979_173_2805_n76), .IN2(
        DP_OP_992_186_8739_n19), .OUT(DP_OP_992_186_8739_n16) );
  NAND2X1 DP_OP_984_178_8739_U34 ( .IN1(n411), .IN2(n407), .OUT(
        DP_OP_984_178_8739_n23) );
  INVX1 DP_OP_987_181_8739_U33 ( .IN(DP_OP_987_181_8739_n23), .OUT(
        DP_OP_987_181_8739_n32) );
  NAND2X1 DP_OP_988_182_8739_U24 ( .IN1(DP_OP_979_173_2805_n76), .IN2(
        DP_OP_988_182_8739_n19), .OUT(DP_OP_988_182_8739_n16) );
  NAND2X1 DP_OP_985_179_8739_U37 ( .IN1(n410), .IN2(DP_OP_985_179_8739_n27), 
        .OUT(DP_OP_985_179_8739_n25) );
  NAND2X1 DP_OP_985_179_8739_U36 ( .IN1(n407), .IN2(DP_OP_985_179_8739_n27), 
        .OUT(DP_OP_985_179_8739_n24) );
  INVX1 DP_OP_980_174_8739_U21 ( .IN(DP_OP_980_174_8739_n15), .OUT(
        DP_OP_980_174_8739_n26) );
  NAND2X1 DP_OP_992_186_8739_U12 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_992_186_8739_n11), .OUT(DP_OP_992_186_8739_n8) );
  INVX1 DP_OP_986_180_8739_U21 ( .IN(DP_OP_986_180_8739_n15), .OUT(
        DP_OP_986_180_8739_n18) );
  INVX1 DP_OP_982_176_8739_U21 ( .IN(DP_OP_982_176_8739_n15), .OUT(
        DP_OP_982_176_8739_n22) );
  NAND2X1 DP_OP_983_177_8739_U30 ( .IN1(n411), .IN2(DP_OP_983_177_8739_n23), 
        .OUT(DP_OP_983_177_8739_n20) );
  INVX1 DP_OP_987_181_8739_U27 ( .IN(DP_OP_987_181_8739_n19), .OUT(
        DP_OP_987_181_8739_n31) );
  INVX1 DP_OP_988_182_8739_U27 ( .IN(DP_OP_988_182_8739_n19), .OUT(
        DP_OP_988_182_8739_n27) );
  NAND2X1 DP_OP_992_186_8739_U18 ( .IN1(DP_OP_979_173_2805_n77), .IN2(
        DP_OP_992_186_8739_n15), .OUT(DP_OP_992_186_8739_n12) );
  INVX1 DP_OP_980_174_8739_U15 ( .IN(DP_OP_980_174_8739_n11), .OUT(
        DP_OP_980_174_8739_n25) );
  INVX1 DP_OP_985_179_8739_U15 ( .IN(DP_OP_985_179_8739_n11), .OUT(
        DP_OP_985_179_8739_n29) );
  INVX1 DP_OP_985_179_8739_U9 ( .IN(DP_OP_985_179_8739_n7), .OUT(
        DP_OP_985_179_8739_n28) );
  INVX1 DP_OP_986_180_8739_U15 ( .IN(DP_OP_986_180_8739_n11), .OUT(
        DP_OP_986_180_8739_n17) );
  INVX1 DP_OP_982_176_8739_U15 ( .IN(DP_OP_982_176_8739_n11), .OUT(
        DP_OP_982_176_8739_n21) );
  INVX1 DP_OP_988_182_8739_U9 ( .IN(DP_OP_988_182_8739_n7), .OUT(
        DP_OP_988_182_8739_n24) );
  INVX4 DP_OP_992_186_8739_U33 ( .IN(DP_OP_992_186_8739_n23), .OUT(
        DP_OP_992_186_8739_n32) );
  NANDX2 DP_OP_992_186_8739_U23 ( .IN1(DP_OP_992_186_8739_n17), .IN2(
        DP_OP_992_186_8739_n16), .OUT(C1_DATA14_3) );
  INVX4 DP_OP_983_177_8739_U33 ( .IN(DP_OP_983_177_8739_n23), .OUT(
        DP_OP_983_177_8739_n32) );
  NANDX2 DP_OP_990_184_2805_U53 ( .IN1(DP_OP_990_184_2805_n22), .IN2(
        DP_OP_990_184_2805_n21), .OUT(C1_DATA12_1) );
  NANDX2 DP_OP_985_179_8739_U35 ( .IN1(DP_OP_985_179_8739_n25), .IN2(
        DP_OP_985_179_8739_n24), .OUT(C1_DATA7_1) );
  INVX4 DP_OP_992_186_8739_U27 ( .IN(DP_OP_992_186_8739_n19), .OUT(
        DP_OP_992_186_8739_n31) );
  INVX4 DP_OP_992_186_8739_U21 ( .IN(DP_OP_992_186_8739_n15), .OUT(
        DP_OP_992_186_8739_n30) );
  NANDX2 DP_OP_992_186_8739_U11 ( .IN1(DP_OP_992_186_8739_n9), .IN2(
        DP_OP_992_186_8739_n8), .OUT(C1_DATA14_5) );
  NANDX2 DP_OP_979_173_2805_U16 ( .IN1(DP_OP_979_173_2805_n10), .IN2(
        DP_OP_979_173_2805_n9), .OUT(C1_DATA1_5) );
  NANDX2 DP_OP_989_183_2805_U16 ( .IN1(DP_OP_989_183_2805_n10), .IN2(
        DP_OP_989_183_2805_n9), .OUT(C1_DATA11_5) );
  NANDX2 DP_OP_991_185_2805_U16 ( .IN1(DP_OP_991_185_2805_n10), .IN2(
        DP_OP_991_185_2805_n9), .OUT(C1_DATA13_5) );
  NANDX2 DP_OP_983_177_8739_U29 ( .IN1(DP_OP_983_177_8739_n21), .IN2(
        DP_OP_983_177_8739_n20), .OUT(C1_DATA5_2) );
  NANDX2 DP_OP_979_173_2805_U44 ( .IN1(DP_OP_979_173_2805_n19), .IN2(
        DP_OP_979_173_2805_n18), .OUT(C1_DATA1_2) );
  NANDX2 DP_OP_979_173_2805_U26 ( .IN1(DP_OP_979_173_2805_n13), .IN2(
        DP_OP_979_173_2805_n12), .OUT(C1_DATA1_4) );
  NANDX2 DP_OP_989_183_2805_U26 ( .IN1(DP_OP_989_183_2805_n13), .IN2(
        DP_OP_989_183_2805_n12), .OUT(C1_DATA11_4) );
  NANDX2 DP_OP_992_186_8739_U17 ( .IN1(DP_OP_992_186_8739_n13), .IN2(
        DP_OP_992_186_8739_n12), .OUT(C1_DATA14_4) );
  INVX4 DP_OP_992_186_8739_U15 ( .IN(DP_OP_992_186_8739_n11), .OUT(
        DP_OP_992_186_8739_n29) );
  NANDX2 DP_OP_985_179_8739_U40 ( .IN1(Final_Exponent_reg[1]), .IN2(
        Final_Exponent_reg[0]), .OUT(DP_OP_985_179_8739_n27) );
  INVX1 DP_OP_984_178_8739_U33 ( .IN(DP_OP_984_178_8739_n23), .OUT(
        DP_OP_984_178_8739_n28) );
  NANDX2 DP_OP_990_184_2805_U17 ( .IN1(n187), .IN2(DP_OP_990_184_2805_n11), 
        .OUT(DP_OP_990_184_2805_n9) );
  NAND2X1 DP_OP_983_177_8739_U31 ( .IN1(n205), .IN2(DP_OP_983_177_8739_n23), 
        .OUT(DP_OP_983_177_8739_n21) );
  NAND2X1 DP_OP_979_173_2805_U46 ( .IN1(DP_OP_979_173_2805_n55), .IN2(
        DP_OP_979_173_2805_n20), .OUT(DP_OP_979_173_2805_n19) );
  NAND2X1 DP_OP_989_183_2805_U28 ( .IN1(DP_OP_989_183_2805_n48), .IN2(
        DP_OP_989_183_2805_n14), .OUT(DP_OP_989_183_2805_n13) );
  INVX1 DP_OP_984_178_8739_U15 ( .IN(DP_OP_984_178_8739_n11), .OUT(
        DP_OP_984_178_8739_n25) );
  INVX1 DP_OP_984_178_8739_U9 ( .IN(DP_OP_984_178_8739_n7), .OUT(
        DP_OP_984_178_8739_n24) );
  NANDX2 DP_OP_992_186_8739_U28 ( .IN1(DP_OP_979_173_2805_n76), .IN2(
        DP_OP_992_186_8739_n32), .OUT(DP_OP_992_186_8739_n19) );
  NAND2X1 DP_OP_992_186_8739_U25 ( .IN1(DP_OP_992_186_8739_n32), .IN2(
        DP_OP_992_186_8739_n19), .OUT(DP_OP_992_186_8739_n17) );
  INVX1 DP_OP_988_182_8739_U33 ( .IN(DP_OP_988_182_8739_n23), .OUT(
        DP_OP_988_182_8739_n28) );
  NAND2X1 DP_OP_988_182_8739_U25 ( .IN1(DP_OP_988_182_8739_n28), .IN2(
        DP_OP_988_182_8739_n19), .OUT(DP_OP_988_182_8739_n17) );
  NAND2X1 DP_OP_989_183_2805_U56 ( .IN1(n201), .IN2(n407), .OUT(
        DP_OP_989_183_2805_n23) );
  NANDX2 DP_OP_992_186_8739_U22 ( .IN1(DP_OP_979_173_2805_n77), .IN2(
        DP_OP_992_186_8739_n31), .OUT(DP_OP_992_186_8739_n15) );
  NANDX2 DP_OP_992_186_8739_U16 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_992_186_8739_n30), .OUT(DP_OP_992_186_8739_n11) );
  NAND2X1 DP_OP_992_186_8739_U19 ( .IN1(DP_OP_992_186_8739_n31), .IN2(
        DP_OP_992_186_8739_n15), .OUT(DP_OP_992_186_8739_n13) );
  NANDX2 DP_OP_992_186_8739_U10 ( .IN1(DP_OP_979_173_2805_n79), .IN2(
        DP_OP_992_186_8739_n29), .OUT(DP_OP_992_186_8739_n7) );
  NANDX2 DP_OP_992_186_8739_U34 ( .IN1(n411), .IN2(n203), .OUT(
        DP_OP_992_186_8739_n23) );
  NANDX2 DP_OP_987_181_8739_U28 ( .IN1(DP_OP_979_173_2805_n76), .IN2(
        DP_OP_987_181_8739_n32), .OUT(DP_OP_987_181_8739_n19) );
  NAND2X1 DP_OP_992_186_8739_U13 ( .IN1(DP_OP_992_186_8739_n30), .IN2(
        DP_OP_992_186_8739_n11), .OUT(DP_OP_992_186_8739_n9) );
  NANDX2 DP_OP_988_182_8739_U28 ( .IN1(DP_OP_979_173_2805_n76), .IN2(
        DP_OP_988_182_8739_n28), .OUT(DP_OP_988_182_8739_n19) );
  NANDX2 DP_OP_983_177_8739_U34 ( .IN1(n411), .IN2(n205), .OUT(
        DP_OP_983_177_8739_n23) );
  NANDX2 DP_OP_990_184_2805_U11 ( .IN1(DP_OP_979_173_2805_n35), .IN2(
        DP_OP_979_173_2805_n45), .OUT(DP_OP_990_184_2805_n34) );
  NAND2X1 DP_OP_982J1_125_6202_U109 ( .IN1(DP_OP_982J1_125_6202_n129), .IN2(
        DP_OP_982J1_125_6202_n113), .OUT(DP_OP_982J1_125_6202_n97) );
  NANDX2 DP_OP_982J1_125_6202_U16 ( .IN1(n200), .IN2(DP_OP_982J1_125_6202_n175), .OUT(DP_OP_982J1_125_6202_n12) );
  NANDX2 DP_OP_982J1_125_6202_U101 ( .IN1(DP_OP_982J1_125_6202_n136), .IN2(
        DP_OP_982J1_125_6202_n180), .OUT(DP_OP_982J1_125_6202_n108) );
  NANDX2 DP_OP_982J1_125_6202_U129 ( .IN1(DP_OP_982J1_125_6202_n131), .IN2(
        DP_OP_982J1_125_6202_n121), .OUT(DP_OP_982J1_125_6202_n99) );
  NANDX2 DP_OP_982J1_125_6202_U29 ( .IN1(DP_OP_982J1_125_6202_n28), .IN2(
        DP_OP_982J1_125_6202_n27), .OUT(N162) );
  NANDX2 DP_OP_982J1_125_6202_U33 ( .IN1(DP_OP_982J1_125_6202_n31), .IN2(
        DP_OP_982J1_125_6202_n4), .OUT(DP_OP_982J1_125_6202_n33) );
  NANDX2 DP_OP_982J1_125_6202_U89 ( .IN1(DP_OP_982J1_125_6202_n127), .IN2(
        DP_OP_982J1_125_6202_n105), .OUT(DP_OP_982J1_125_6202_n95) );
  NANDX2 DP_OP_982J1_125_6202_U98 ( .IN1(DP_OP_982J1_125_6202_n128), .IN2(
        DP_OP_982J1_125_6202_n108), .OUT(DP_OP_982J1_125_6202_n96) );
  NANDX2 DP_OP_982J1_125_6202_U132 ( .IN1(DP_OP_982J1_125_6202_n139), .IN2(
        DP_OP_982J1_125_6202_n177), .OUT(DP_OP_982J1_125_6202_n121) );
  NANDX2 DP_OP_982J1_125_6202_U133 ( .IN1(DP_OP_982J1_125_6202_n90), .IN2(
        DP_OP_982J1_125_6202_n89), .OUT(N419) );
  NANDX2 DP_OP_982J1_125_6202_U138 ( .IN1(DP_OP_982J1_125_6202_n132), .IN2(
        DP_OP_982J1_125_6202_n124), .OUT(DP_OP_982J1_125_6202_n100) );
  NOR2X1 DP_OP_982J1_125_6202_U142 ( .IN1(DP_OP_982J1_125_6202_n35), .IN2(
        DP_OP_982J1_125_6202_n34), .OUT(N418) );
  NOR2X1 DP_OP_982J1_125_6202_U140 ( .IN1(Datain2[8]), .IN2(n272), .OUT(
        DP_OP_982J1_125_6202_n123) );
  OAI21 DP_OP_982J1_125_6202_U137 ( .IN1(n204), .IN2(DP_OP_982J1_125_6202_n123), .IN3(DP_OP_982J1_125_6202_n124), .OUT(DP_OP_982J1_125_6202_n122) );
  NOR2X1 DP_OP_982J1_125_6202_U131 ( .IN1(DP_OP_982J1_125_6202_n177), .IN2(
        DP_OP_982J1_125_6202_n139), .OUT(DP_OP_982J1_125_6202_n120) );
  NAND2X1 DP_OP_982J1_125_6202_U112 ( .IN1(DP_OP_982J1_125_6202_n137), .IN2(
        Datain2[11]), .OUT(DP_OP_982J1_125_6202_n113) );
  NOR2X1 DP_OP_982J1_125_6202_U111 ( .IN1(Datain2[11]), .IN2(
        DP_OP_982J1_125_6202_n137), .OUT(DP_OP_982J1_125_6202_n112) );
  NOR2X1 DP_OP_982J1_125_6202_U100 ( .IN1(DP_OP_982J1_125_6202_n180), .IN2(
        DP_OP_982J1_125_6202_n136), .OUT(DP_OP_982J1_125_6202_n107) );
  NAND2X1 DP_OP_982J1_125_6202_U92 ( .IN1(DP_OP_982J1_125_6202_n135), .IN2(
        DP_OP_982J1_125_6202_n181), .OUT(DP_OP_982J1_125_6202_n105) );
  NOR2X1 DP_OP_982J1_125_6202_U91 ( .IN1(DP_OP_982J1_125_6202_n181), .IN2(
        DP_OP_982J1_125_6202_n135), .OUT(DP_OP_982J1_125_6202_n104) );
  NOR2X1 DP_OP_982J1_125_6202_U82 ( .IN1(DP_OP_982J1_125_6202_n75), .IN2(
        DP_OP_982J1_125_6202_n74), .OUT(N424) );
  FULLADD DP_OP_982J1_125_6202_U66 ( .A(n272), .B(Datain2[8]), .CIN(
        DP_OP_982J1_125_6202_n63), .COUT(DP_OP_982J1_125_6202_n62), .SUM(N156)
         );
  FULLADD DP_OP_982J1_125_6202_U65 ( .A(DP_OP_982J1_125_6202_n139), .B(
        DP_OP_982J1_125_6202_n177), .CIN(DP_OP_982J1_125_6202_n62), .COUT(
        DP_OP_982J1_125_6202_n61), .SUM(N157) );
  NOR2X1 DP_OP_982J1_125_6202_U45 ( .IN1(DP_OP_982J1_125_6202_n16), .IN2(
        DP_OP_982J1_125_6202_n15), .OUT(DP_OP_982J1_125_6202_n44) );
  FULLADD DP_OP_982J1_125_6202_U38 ( .A(DP_OP_981J1_124_6202_n140), .B(n272), 
        .CIN(n226), .COUT(DP_OP_982J1_125_6202_n38), .SUM(N160) );
  FULLADD DP_OP_982J1_125_6202_U37 ( .A(DP_OP_982J1_125_6202_n24), .B(
        DP_OP_982J1_125_6202_n139), .CIN(DP_OP_982J1_125_6202_n38), .COUT(
        DP_OP_982J1_125_6202_n37), .SUM(N161) );
  NOR2X1 DP_OP_982J1_125_6202_U21 ( .IN1(DP_OP_982J1_125_6202_n20), .IN2(
        DP_OP_982J1_125_6202_n45), .OUT(DP_OP_982J1_125_6202_n24) );
  NAND2X1 DP_OP_982J1_125_6202_U13 ( .IN1(DP_OP_982J1_125_6202_n66), .IN2(
        DP_OP_982J1_125_6202_n12), .OUT(DP_OP_982J1_125_6202_n8) );
  FULLADD DP_OP_982J1_125_6202_U10 ( .A(DP_OP_981J1_124_6202_n140), .B(n272), 
        .CIN(DP_OP_982J1_125_6202_n63), .COUT(DP_OP_982J1_125_6202_n10), .SUM(
        N164) );
  FULLADD DP_OP_982J1_125_6202_U9 ( .A(n191), .B(DP_OP_982J1_125_6202_n139), 
        .CIN(DP_OP_982J1_125_6202_n10), .COUT(DP_OP_982J1_125_6202_n9), .SUM(
        N165) );
  NANDX2 DP_OP_981J1_124_6202_U113 ( .IN1(DP_OP_981J1_124_6202_n84), .IN2(
        DP_OP_981J1_124_6202_n83), .OUT(N365) );
  NANDX2 DP_OP_981J1_124_6202_U132 ( .IN1(n220), .IN2(Datain1[9]), .OUT(
        DP_OP_981J1_124_6202_n121) );
  NAND2X1 DP_OP_981J1_124_6202_U138 ( .IN1(n241), .IN2(
        DP_OP_981J1_124_6202_n124), .OUT(DP_OP_981J1_124_6202_n100) );
  NAND2X1 DP_OP_981J1_124_6202_U118 ( .IN1(DP_OP_982J1_125_6202_n58), .IN2(
        DP_OP_982J1_125_6202_n130), .OUT(DP_OP_981J1_124_6202_n98) );
  NANDX2 DP_OP_981J1_124_6202_U33 ( .IN1(DP_OP_981J1_124_6202_n31), .IN2(
        DP_OP_981J1_124_6202_n4), .OUT(DP_OP_981J1_124_6202_n33) );
  NANDX2 DP_OP_981J1_124_6202_U133 ( .IN1(DP_OP_981J1_124_6202_n90), .IN2(
        DP_OP_981J1_124_6202_n89), .OUT(N363) );
  NANDX2 DP_OP_981J1_124_6202_U89 ( .IN1(DP_OP_981J1_124_6202_n127), .IN2(
        DP_OP_981J1_124_6202_n105), .OUT(DP_OP_981J1_124_6202_n95) );
  NANDX2 DP_OP_981J1_124_6202_U98 ( .IN1(n237), .IN2(DP_OP_981J1_124_6202_n108), .OUT(DP_OP_981J1_124_6202_n96) );
  NOR2X1 DP_OP_981J1_124_6202_U140 ( .IN1(Datain1[8]), .IN2(
        DP_OP_981J1_124_6202_n140), .OUT(DP_OP_981J1_124_6202_n123) );
  NOR2X1 DP_OP_981J1_124_6202_U131 ( .IN1(Datain1[9]), .IN2(n220), .OUT(
        DP_OP_981J1_124_6202_n120) );
  NAND2X1 DP_OP_981J1_124_6202_U112 ( .IN1(DP_OP_981J1_124_6202_n137), .IN2(
        Datain1[11]), .OUT(DP_OP_981J1_124_6202_n113) );
  NOR2X1 DP_OP_981J1_124_6202_U111 ( .IN1(Datain1[11]), .IN2(
        DP_OP_981J1_124_6202_n137), .OUT(DP_OP_981J1_124_6202_n112) );
  NAND2X1 DP_OP_981J1_124_6202_U109 ( .IN1(DP_OP_981J1_124_6202_n129), .IN2(
        DP_OP_981J1_124_6202_n113), .OUT(DP_OP_981J1_124_6202_n97) );
  NAND2X1 DP_OP_981J1_124_6202_U101 ( .IN1(n206), .IN2(Datain1[12]), .OUT(
        DP_OP_981J1_124_6202_n108) );
  NOR2X1 DP_OP_981J1_124_6202_U100 ( .IN1(Datain1[12]), .IN2(n206), .OUT(
        DP_OP_981J1_124_6202_n107) );
  NAND2X1 DP_OP_981J1_124_6202_U92 ( .IN1(DP_OP_981J1_124_6202_n135), .IN2(
        Datain1[13]), .OUT(DP_OP_981J1_124_6202_n105) );
  NOR2X1 DP_OP_981J1_124_6202_U91 ( .IN1(Datain1[13]), .IN2(
        DP_OP_981J1_124_6202_n135), .OUT(DP_OP_981J1_124_6202_n104) );
  FULLADD DP_OP_981J1_124_6202_U66 ( .A(DP_OP_981J1_124_6202_n140), .B(
        Datain1[8]), .CIN(n204), .COUT(DP_OP_981J1_124_6202_n62), .SUM(N144)
         );
  FULLADD DP_OP_981J1_124_6202_U65 ( .A(n220), .B(Datain1[9]), .CIN(
        DP_OP_981J1_124_6202_n62), .COUT(DP_OP_981J1_124_6202_n61), .SUM(N145)
         );
  NOR2X1 DP_OP_981J1_124_6202_U45 ( .IN1(DP_OP_981J1_124_6202_n16), .IN2(
        DP_OP_981J1_124_6202_n15), .OUT(DP_OP_981J1_124_6202_n44) );
  FULLADD DP_OP_981J1_124_6202_U38 ( .A(n272), .B(DP_OP_981J1_124_6202_n140), 
        .CIN(n250), .COUT(DP_OP_981J1_124_6202_n38), .SUM(N148) );
  FULLADD DP_OP_981J1_124_6202_U37 ( .A(n190), .B(n220), .CIN(
        DP_OP_981J1_124_6202_n38), .COUT(DP_OP_981J1_124_6202_n37), .SUM(N149)
         );
  NOR2X1 DP_OP_981J1_124_6202_U21 ( .IN1(DP_OP_981J1_124_6202_n20), .IN2(
        DP_OP_981J1_124_6202_n45), .OUT(DP_OP_981J1_124_6202_n24) );
  NAND2X1 DP_OP_981J1_124_6202_U13 ( .IN1(n250), .IN2(DP_OP_982J1_125_6202_n66), .OUT(DP_OP_981J1_124_6202_n8) );
  FULLADD DP_OP_981J1_124_6202_U10 ( .A(n272), .B(DP_OP_981J1_124_6202_n140), 
        .CIN(n204), .COUT(DP_OP_981J1_124_6202_n10), .SUM(N152) );
  FULLADD DP_OP_981J1_124_6202_U9 ( .A(DP_OP_981J1_124_6202_n24), .B(n220), 
        .CIN(DP_OP_981J1_124_6202_n10), .COUT(DP_OP_981J1_124_6202_n9), .SUM(
        N153) );
  NANDX2 DP_OP_982J1_125_6202_U141 ( .IN1(n272), .IN2(Datain2[8]), .OUT(
        DP_OP_982J1_125_6202_n124) );
  NANDX2 DP_OP_981J1_124_6202_U129 ( .IN1(DP_OP_981J1_124_6202_n131), .IN2(
        DP_OP_981J1_124_6202_n121), .OUT(DP_OP_981J1_124_6202_n99) );
  NAND2X1 DP_OP_992_186_8739_U35 ( .IN1(DP_OP_985_179_8739_n25), .IN2(
        DP_OP_985_179_8739_n24), .OUT(C1_DATA14_1) );
  NAND2X1 DP_OP_988_182_8739_U23 ( .IN1(DP_OP_988_182_8739_n17), .IN2(
        DP_OP_988_182_8739_n16), .OUT(C1_DATA10_3) );
  NAND2X1 DP_OP_990_184_2805_U54 ( .IN1(n407), .IN2(DP_OP_990_184_2805_n23), 
        .OUT(DP_OP_990_184_2805_n21) );
  NAND2X1 DP_OP_990_184_2805_U5 ( .IN1(DP_OP_990_184_2805_n2), .IN2(
        DP_OP_979_173_2805_n80), .OUT(DP_OP_990_184_2805_n5) );
  NAND2X1 DP_OP_990_184_2805_U29 ( .IN1(DP_OP_990_184_2805_n48), .IN2(
        DP_OP_979_173_2805_n77), .OUT(DP_OP_990_184_2805_n14) );
  NAND2X1 DP_OP_989_183_2805_U29 ( .IN1(DP_OP_989_183_2805_n48), .IN2(
        DP_OP_979_173_2805_n77), .OUT(DP_OP_989_183_2805_n14) );
  NAND2X1 DP_OP_991_185_2805_U29 ( .IN1(DP_OP_991_185_2805_n48), .IN2(
        DP_OP_979_173_2805_n77), .OUT(DP_OP_991_185_2805_n14) );
  NAND2X1 DP_OP_989_183_2805_U9 ( .IN1(DP_OP_989_183_2805_n38), .IN2(
        DP_OP_979_173_2805_n79), .OUT(DP_OP_989_183_2805_n8) );
  NAND2X1 DP_OP_989_183_2805_U5 ( .IN1(DP_OP_989_183_2805_n2), .IN2(
        DP_OP_979_173_2805_n80), .OUT(DP_OP_989_183_2805_n5) );
  NAND2X1 DP_OP_991_185_2805_U5 ( .IN1(DP_OP_991_185_2805_n2), .IN2(
        DP_OP_979_173_2805_n80), .OUT(DP_OP_991_185_2805_n5) );
  NAND2X1 DP_OP_990_184_2805_U16 ( .IN1(DP_OP_990_184_2805_n10), .IN2(
        DP_OP_990_184_2805_n9), .OUT(C1_DATA12_5) );
  NAND2X1 DP_OP_991_185_2805_U19 ( .IN1(DP_OP_991_185_2805_n43), .IN2(
        DP_OP_979_173_2805_n78), .OUT(DP_OP_991_185_2805_n11) );
  NAND2X1 DP_OP_989_183_2805_U19 ( .IN1(DP_OP_989_183_2805_n43), .IN2(
        DP_OP_979_173_2805_n78), .OUT(DP_OP_989_183_2805_n11) );
  NAND2X1 DP_OP_991_185_2805_U3 ( .IN1(DP_OP_979_173_2805_n80), .IN2(
        DP_OP_991_185_2805_n5), .OUT(DP_OP_991_185_2805_n3) );
  NAND2X1 DP_OP_989_183_2805_U3 ( .IN1(DP_OP_979_173_2805_n80), .IN2(
        DP_OP_989_183_2805_n5), .OUT(DP_OP_989_183_2805_n3) );
  NAND2X1 DP_OP_989_183_2805_U27 ( .IN1(DP_OP_979_173_2805_n77), .IN2(
        DP_OP_989_183_2805_n14), .OUT(DP_OP_989_183_2805_n12) );
  NAND2X1 DP_OP_989_183_2805_U17 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_989_183_2805_n11), .OUT(DP_OP_989_183_2805_n9) );
  NAND2X1 DP_OP_991_185_2805_U17 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_991_185_2805_n11), .OUT(DP_OP_991_185_2805_n9) );
  NAND2X1 DP_OP_979_173_2805_U19 ( .IN1(DP_OP_979_173_2805_n43), .IN2(
        DP_OP_979_173_2805_n78), .OUT(DP_OP_979_173_2805_n11) );
  NAND2X1 DP_OP_979_173_2805_U27 ( .IN1(DP_OP_979_173_2805_n77), .IN2(
        DP_OP_979_173_2805_n14), .OUT(DP_OP_979_173_2805_n12) );
  NAND2X1 DP_OP_979_173_2805_U17 ( .IN1(DP_OP_979_173_2805_n78), .IN2(
        DP_OP_979_173_2805_n11), .OUT(DP_OP_979_173_2805_n9) );
  INVX1 DP_OP_979_173_2805_U31 ( .IN(DP_OP_979_173_2805_n45), .OUT(
        DP_OP_979_173_2805_n44) );
  NANDX2 DP_OP_982J1_125_6202_U118 ( .IN1(DP_OP_982J1_125_6202_n130), .IN2(
        DP_OP_982J1_125_6202_n58), .OUT(DP_OP_982J1_125_6202_n98) );
  BUF4X U3 ( .IN(Datain2[9]), .OUT(DP_OP_982J1_125_6202_n177) );
  INVX4 U4 ( .IN(n292), .OUT(n410) );
  BUF4X U5 ( .IN(N418), .OUT(n202) );
  NOR2X1 U6 ( .IN1(n1017), .IN2(n393), .OUT(n1) );
  NAND3X1 U7 ( .IN1(n946), .IN2(n948), .IN3(n1), .OUT(n994) );
  INVX1 U8 ( .IN(DP_OP_979_173_2805_n58), .OUT(n2) );
  MUX2X1 U9 ( .IN1(DP_OP_979_173_2805_n58), .IN2(n2), .S(n407), .OUT(n3) );
  NAND2X1 U10 ( .IN1(n1197), .IN2(n3), .OUT(n1145) );
  INVX1 U11 ( .IN(DP_OP_987_181_8739_n7), .OUT(n4) );
  MUX2X1 U12 ( .IN1(DP_OP_987_181_8739_n7), .IN2(n4), .S(
        DP_OP_979_173_2805_n80), .OUT(C1_DATA9_7) );
  INVX1 U13 ( .IN(DP_OP_979_173_2805_n79), .OUT(n5) );
  INVX1 U14 ( .IN(DP_OP_983_177_8739_n29), .OUT(n6) );
  OAI21 U15 ( .IN1(n5), .IN2(n6), .IN3(DP_OP_983_177_8739_n28), .OUT(
        C1_DATA5_6) );
  INVX1 U16 ( .IN(DP_OP_989_183_2805_n1), .OUT(n7) );
  INVX1 U17 ( .IN(DP_OP_979_173_2805_n76), .OUT(n8) );
  AOI22 U18 ( .IN1(DP_OP_979_173_2805_n76), .IN2(n7), .IN3(
        DP_OP_989_183_2805_n1), .IN4(n8), .OUT(C1_DATA11_3) );
  INVX1 U19 ( .IN(n411), .OUT(n9) );
  INVX1 U20 ( .IN(DP_OP_990_184_2805_n58), .OUT(n10) );
  NOR2X1 U21 ( .IN1(n407), .IN2(n10), .OUT(n11) );
  MUX2X1 U22 ( .IN1(n411), .IN2(n9), .S(n11), .OUT(C1_DATA12_2) );
  INVX1 U23 ( .IN(N165), .OUT(n12) );
  NOR2X1 U24 ( .IN1(N164), .IN2(n12), .OUT(n716) );
  AOI22 U25 ( .IN1(n1179), .IN2(DP_OP_979_173_2805_n76), .IN3(n1564), .IN4(
        Datain2[10]), .OUT(n13) );
  NAND2X1 U26 ( .IN1(n197), .IN2(Datain1[10]), .OUT(n14) );
  NAND2X1 U27 ( .IN1(n13), .IN2(n14), .OUT(n184) );
  OAI21 U28 ( .IN1(Datain1[14]), .IN2(n209), .IN3(n436), .OUT(n15) );
  INVX1 U29 ( .IN(n15), .OUT(DP_OP_982J1_125_6202_n73) );
  INVX1 U30 ( .IN(DP_OP_979_173_2805_n80), .OUT(n16) );
  MUX2X1 U31 ( .IN1(n16), .IN2(DP_OP_979_173_2805_n80), .S(
        DP_OP_984_178_8739_n24), .OUT(C1_DATA6_7) );
  AOI21 U32 ( .IN1(n1210), .IN2(n945), .IN3(n944), .OUT(n17) );
  INVX1 U33 ( .IN(n17), .OUT(n18) );
  NOR2X1 U34 ( .IN1(n998), .IN2(n18), .OUT(n1040) );
  AOI21 U35 ( .IN1(DP_OP_979_173_2805_n79), .IN2(DP_OP_988_182_8739_n25), 
        .IN3(DP_OP_988_182_8739_n7), .OUT(n19) );
  INVX1 U36 ( .IN(n19), .OUT(C1_DATA10_6) );
  INVX1 U37 ( .IN(DP_OP_979_173_2805_n76), .OUT(n20) );
  MUX2X1 U38 ( .IN1(n20), .IN2(DP_OP_979_173_2805_n76), .S(
        DP_OP_989_183_2805_n1), .OUT(C1_DATA13_3) );
  INVX1 U39 ( .IN(n411), .OUT(n21) );
  MUX2X1 U40 ( .IN1(n411), .IN2(n21), .S(DP_OP_989_183_2805_n55), .OUT(
        C1_DATA11_2) );
  INVX1 U41 ( .IN(N149), .OUT(n22) );
  NOR2X1 U42 ( .IN1(N148), .IN2(n22), .OUT(n771) );
  INVX1 U43 ( .IN(DP_OP_980_174_8739_n7), .OUT(n23) );
  MUX2X1 U44 ( .IN1(DP_OP_980_174_8739_n7), .IN2(n23), .S(
        DP_OP_979_173_2805_n80), .OUT(C1_DATA2_7) );
  AOI21 U45 ( .IN1(n185), .IN2(DP_OP_981_175_8739_n32), .IN3(n369), .OUT(n24)
         );
  INVX1 U46 ( .IN(n24), .OUT(C1_DATA3_3) );
  NAND2X1 U47 ( .IN1(n410), .IN2(n921), .OUT(n25) );
  OAI21 U48 ( .IN1(DP_OP_979_173_2805_n58), .IN2(n26), .IN3(n1197), .OUT(n1111) );
  INVX1 U49 ( .IN(n25), .OUT(n26) );
  INVX1 U50 ( .IN(DP_OP_981J1_124_6202_n73), .OUT(n27) );
  MUX2X1 U51 ( .IN1(DP_OP_981J1_124_6202_n73), .IN2(n27), .S(n231), .OUT(N369)
         );
  INVX1 U52 ( .IN(DP_OP_979_173_2805_n80), .OUT(n28) );
  INVX1 U53 ( .IN(DP_OP_982_176_8739_n7), .OUT(n29) );
  AOI22 U54 ( .IN1(DP_OP_982_176_8739_n7), .IN2(DP_OP_979_173_2805_n80), .IN3(
        n28), .IN4(n29), .OUT(C1_DATA4_7) );
  AOI21 U55 ( .IN1(DP_OP_979_173_2805_n79), .IN2(DP_OP_987_181_8739_n29), 
        .IN3(DP_OP_987_181_8739_n7), .OUT(n30) );
  INVX1 U56 ( .IN(n30), .OUT(C1_DATA9_6) );
  INVX1 U57 ( .IN(n890), .OUT(n31) );
  NAND3X1 U58 ( .IN1(n874), .IN2(n591), .IN3(n31), .OUT(n642) );
  INVX1 U59 ( .IN(N157), .OUT(n32) );
  NOR2X1 U60 ( .IN1(N156), .IN2(n32), .OUT(n816) );
  AOI21 U61 ( .IN1(DP_OP_979_173_2805_n79), .IN2(DP_OP_980_174_8739_n25), 
        .IN3(DP_OP_980_174_8739_n7), .OUT(n33) );
  INVX1 U62 ( .IN(n33), .OUT(n34) );
  INVX1 U63 ( .IN(C1_DATA7_6), .OUT(n35) );
  OAI21 U64 ( .IN1(n1184), .IN2(n35), .IN3(n1155), .OUT(n36) );
  AOI21 U65 ( .IN1(n1186), .IN2(n34), .IN3(n36), .OUT(n1162) );
  INVX1 U66 ( .IN(DP_OP_981J1_124_6202_n33), .OUT(n37) );
  MUX2X1 U67 ( .IN1(DP_OP_981J1_124_6202_n33), .IN2(n37), .S(
        DP_OP_981J1_124_6202_n9), .OUT(N154) );
  AOI22 U68 ( .IN1(n306), .IN2(Op1_Sign_reg), .IN3(n305), .IN4(Op2_Sign_reg), 
        .OUT(n38) );
  INVX4 U69 ( .IN(n38), .OUT(n1556) );
  OAI21 U70 ( .IN1(n410), .IN2(n407), .IN3(DP_OP_985_179_8739_n27), .OUT(n39)
         );
  INVX1 U71 ( .IN(n39), .OUT(C1_DATA3_1) );
  AOI21 U72 ( .IN1(n185), .IN2(DP_OP_992_186_8739_n32), .IN3(
        DP_OP_985_179_8739_n19), .OUT(n1049) );
  NOR2X1 U73 ( .IN1(DP_OP_988_182_8739_n13), .IN2(DP_OP_988_182_8739_n12), 
        .OUT(n40) );
  AOI21 U74 ( .IN1(DP_OP_979_173_2805_n77), .IN2(DP_OP_983_177_8739_n31), 
        .IN3(DP_OP_983_177_8739_n15), .OUT(n41) );
  INVX1 U75 ( .IN(n41), .OUT(n42) );
  AOI22 U76 ( .IN1(n1192), .IN2(n40), .IN3(n1191), .IN4(n42), .OUT(n1169) );
  INVX1 U77 ( .IN(n411), .OUT(n43) );
  MUX2X1 U78 ( .IN1(n411), .IN2(n43), .S(DP_OP_989_183_2805_n55), .OUT(
        C1_DATA13_2) );
  NAND3X1 U79 ( .IN1(n425), .IN2(n615), .IN3(n423), .OUT(n891) );
  INVX1 U80 ( .IN(DP_OP_979_173_2805_n79), .OUT(n44) );
  NOR2X1 U81 ( .IN1(DP_OP_990_184_2805_n51), .IN2(DP_OP_979_173_2805_n39), 
        .OUT(n45) );
  MUX2X1 U82 ( .IN1(DP_OP_979_173_2805_n79), .IN2(n44), .S(n45), .OUT(n46) );
  NAND2X1 U83 ( .IN1(n1272), .IN2(n46), .OUT(n328) );
  NAND3X1 U84 ( .IN1(DP_OP_982J1_125_6202_n135), .IN2(
        DP_OP_982J1_125_6202_n136), .IN3(n1615), .OUT(n47) );
  NAND3X1 U85 ( .IN1(n259), .IN2(n200), .IN3(n272), .OUT(n48) );
  NOR2X1 U86 ( .IN1(n47), .IN2(n48), .OUT(n49) );
  NAND3X1 U87 ( .IN1(DP_OP_982J1_125_6202_n137), .IN2(
        DP_OP_982J1_125_6202_n139), .IN3(n49), .OUT(n1621) );
  AOI22 U88 ( .IN1(Datain2[8]), .IN2(n768), .IN3(n767), .IN4(
        DP_OP_982J1_125_6202_n182), .OUT(n50) );
  OAI21 U89 ( .IN1(n1570), .IN2(n770), .IN3(n769), .OUT(n51) );
  AOI21 U90 ( .IN1(DP_OP_982J1_125_6202_n180), .IN2(n771), .IN3(n51), .OUT(n52) );
  OAI21 U91 ( .IN1(DP_OP_981J1_124_6202_n137), .IN2(n770), .IN3(N147), .OUT(
        n53) );
  AOI21 U92 ( .IN1(DP_OP_982J1_125_6202_n181), .IN2(n771), .IN3(n53), .OUT(n54) );
  AOI22 U93 ( .IN1(DP_OP_982J1_125_6202_n177), .IN2(n768), .IN3(n767), .IN4(
        Datain2[15]), .OUT(n55) );
  AOI22 U94 ( .IN1(n50), .IN2(n52), .IN3(n54), .IN4(n55), .OUT(n56) );
  INVX1 U95 ( .IN(n56), .OUT(n327) );
  NOR2X1 U96 ( .IN1(n1185), .IN2(n1196), .OUT(n57) );
  AOI22 U97 ( .IN1(n1186), .IN2(C1_DATA2_7), .IN3(n1197), .IN4(C1_DATA1_7), 
        .OUT(n58) );
  NAND2X1 U98 ( .IN1(n57), .IN2(n58), .OUT(n348) );
  AOI22 U99 ( .IN1(n1482), .IN2(n1499), .IN3(n1483), .IN4(
        Final_Mantissa_reg[10]), .OUT(n59) );
  OAI21 U100 ( .IN1(n1485), .IN2(n1484), .IN3(n59), .OUT(n60) );
  AOI22 U101 ( .IN1(Debug_reg[0]), .IN2(n1535), .IN3(n1534), .IN4(n60), .OUT(
        n61) );
  INVX1 U102 ( .IN(n61), .OUT(n109) );
  AOI21 U103 ( .IN1(DP_OP_979_173_2805_n78), .IN2(DP_OP_986_180_8739_n18), 
        .IN3(DP_OP_986_180_8739_n11), .OUT(n62) );
  INVX1 U104 ( .IN(n62), .OUT(C1_DATA8_5) );
  OAI21 U105 ( .IN1(DP_OP_991_185_2805_n48), .IN2(DP_OP_979_173_2805_n77), 
        .IN3(DP_OP_991_185_2805_n14), .OUT(n63) );
  INVX1 U106 ( .IN(n63), .OUT(C1_DATA13_4) );
  OAI21 U107 ( .IN1(n203), .IN2(n411), .IN3(DP_OP_992_186_8739_n23), .OUT(n64)
         );
  INVX1 U108 ( .IN(n64), .OUT(C1_DATA14_2) );
  INVX1 U109 ( .IN(DP_OP_982J1_125_6202_n97), .OUT(n65) );
  OAI21 U110 ( .IN1(DP_OP_982J1_125_6202_n117), .IN2(n273), .IN3(
        DP_OP_982J1_125_6202_n58), .OUT(n66) );
  MUX2X1 U111 ( .IN1(n65), .IN2(DP_OP_982J1_125_6202_n97), .S(n66), .OUT(N422)
         );
  AOI21 U112 ( .IN1(DP_OP_979_173_2805_n77), .IN2(DP_OP_982_176_8739_n23), 
        .IN3(DP_OP_982_176_8739_n15), .OUT(n67) );
  INVX1 U113 ( .IN(n67), .OUT(n68) );
  INVX1 U114 ( .IN(DP_OP_987_181_8739_n15), .OUT(n69) );
  INVX1 U115 ( .IN(DP_OP_979_173_2805_n77), .OUT(n70) );
  AOI21 U116 ( .IN1(n69), .IN2(n70), .IN3(DP_OP_987_181_8739_n13), .OUT(n71)
         );
  AOI22 U117 ( .IN1(n1190), .IN2(n68), .IN3(n1189), .IN4(n71), .OUT(n1170) );
  NAND3X1 U118 ( .IN1(DP_OP_979_173_2805_n77), .IN2(DP_OP_979_173_2805_n78), 
        .IN3(DP_OP_979_173_2805_n80), .OUT(n72) );
  NAND3X1 U119 ( .IN1(n411), .IN2(n407), .IN3(DP_OP_979_173_2805_n79), .OUT(
        n74) );
  NOR2X1 U120 ( .IN1(n72), .IN2(n74), .OUT(n75) );
  NAND3X1 U121 ( .IN1(n410), .IN2(DP_OP_979_173_2805_n76), .IN3(n75), .OUT(
        n977) );
  INVX1 U122 ( .IN(N145), .OUT(n76) );
  NOR2X1 U123 ( .IN1(N144), .IN2(n76), .OUT(n841) );
  INVX1 U124 ( .IN(DP_OP_979_173_2805_n80), .OUT(n77) );
  MUX2X1 U125 ( .IN1(n77), .IN2(DP_OP_979_173_2805_n80), .S(
        DP_OP_992_186_8739_n7), .OUT(C1_DATA14_7) );
  INVX1 U126 ( .IN(DP_OP_986_180_8739_n7), .OUT(n78) );
  MUX2X1 U127 ( .IN1(DP_OP_986_180_8739_n7), .IN2(n78), .S(
        DP_OP_979_173_2805_n80), .OUT(C1_DATA8_7) );
  INVX1 U128 ( .IN(DP_OP_979_173_2805_n80), .OUT(n79) );
  NOR2X1 U129 ( .IN1(DP_OP_990_184_2805_n34), .IN2(DP_OP_979_173_2805_n1), 
        .OUT(n80) );
  MUX2X1 U130 ( .IN1(DP_OP_979_173_2805_n80), .IN2(n79), .S(n80), .OUT(
        C1_DATA1_7) );
  NAND3X1 U131 ( .IN1(n1487), .IN2(n1219), .IN3(n928), .OUT(n81) );
  INVX1 U132 ( .IN(n81), .OUT(n82) );
  NAND3X1 U133 ( .IN1(n936), .IN2(n1493), .IN3(n82), .OUT(n1482) );
  INVX1 U134 ( .IN(n1479), .OUT(n83) );
  NAND3X1 U135 ( .IN1(add_x_35_A_2_), .IN2(add_x_35_A_3_), .IN3(n83), .OUT(
        n1551) );
  INVX1 U136 ( .IN(DP_OP_982J1_125_6202_n33), .OUT(n84) );
  MUX2X1 U137 ( .IN1(DP_OP_982J1_125_6202_n33), .IN2(n84), .S(
        DP_OP_982J1_125_6202_n9), .OUT(N166) );
  AOI22 U138 ( .IN1(n768), .IN2(Datain2[1]), .IN3(n771), .IN4(Datain2[5]), 
        .OUT(n85) );
  OAI21 U139 ( .IN1(n86), .IN2(n87), .IN3(n85), .OUT(n88) );
  AOI22 U140 ( .IN1(n768), .IN2(Datain2[0]), .IN3(n771), .IN4(Datain2[4]), 
        .OUT(n89) );
  AOI21 U141 ( .IN1(n767), .IN2(Datain2[6]), .IN3(n766), .OUT(n90) );
  NAND2X1 U142 ( .IN1(n89), .IN2(n90), .OUT(n91) );
  OAI21 U143 ( .IN1(n764), .IN2(n88), .IN3(n91), .OUT(n326) );
  INVX1 U144 ( .IN(Datain2[7]), .OUT(n86) );
  INVX1 U145 ( .IN(n767), .OUT(n87) );
  NAND3X1 U146 ( .IN1(n1160), .IN2(n1161), .IN3(n1163), .OUT(n92) );
  NAND2X1 U147 ( .IN1(n328), .IN2(n1162), .OUT(n93) );
  OAI21 U148 ( .IN1(n92), .IN2(n93), .IN3(n1534), .OUT(n94) );
  NAND3X1 U149 ( .IN1(n1165), .IN2(n1164), .IN3(n94), .OUT(n1100) );
  INVX1 U150 ( .IN(DP_OP_982J1_125_6202_n105), .OUT(n95) );
  AOI21 U151 ( .IN1(DP_OP_982J1_125_6202_n127), .IN2(n285), .IN3(n95), .OUT(
        n289) );
  INVX1 U152 ( .IN(DP_OP_985_179_8739_n30), .OUT(n96) );
  AOI21 U153 ( .IN1(DP_OP_985_179_8739_n31), .IN2(DP_OP_979_173_2805_n77), 
        .IN3(n96), .OUT(n1167) );
  OAI21 U154 ( .IN1(n407), .IN2(n411), .IN3(DP_OP_984_178_8739_n23), .OUT(n97)
         );
  INVX1 U155 ( .IN(n97), .OUT(C1_DATA6_2) );
  AOI21 U156 ( .IN1(n411), .IN2(n203), .IN3(DP_OP_981_175_8739_n23), .OUT(n98)
         );
  INVX1 U157 ( .IN(n98), .OUT(C1_DATA3_2) );
  INVX1 U158 ( .IN(n1615), .OUT(n99) );
  MUX2X1 U159 ( .IN1(n1615), .IN2(n99), .S(DP_OP_982J1_125_6202_n182), .OUT(
        DP_OP_981J1_124_6202_n73) );
  AOI21 U160 ( .IN1(n411), .IN2(n407), .IN3(n210), .OUT(n100) );
  INVX1 U161 ( .IN(n100), .OUT(C1_DATA2_2) );
  INVX1 U162 ( .IN(DP_OP_981J1_124_6202_n95), .OUT(n101) );
  MUX2X1 U163 ( .IN1(n101), .IN2(DP_OP_981J1_124_6202_n95), .S(
        DP_OP_981J1_124_6202_n106), .OUT(N368) );
  NAND3X1 U164 ( .IN1(n438), .IN2(n345), .IN3(n1621), .OUT(n1316) );
  NAND3X1 U165 ( .IN1(n937), .IN2(n942), .IN3(n1003), .OUT(n1251) );
  AOI21 U166 ( .IN1(DP_OP_979_173_2805_n79), .IN2(DP_OP_985_179_8739_n29), 
        .IN3(DP_OP_985_179_8739_n7), .OUT(n102) );
  INVX1 U167 ( .IN(n102), .OUT(C1_DATA7_6) );
  AOI21 U168 ( .IN1(DP_OP_979_173_2805_n79), .IN2(DP_OP_982_176_8739_n21), 
        .IN3(DP_OP_982_176_8739_n7), .OUT(n104) );
  INVX1 U169 ( .IN(n104), .OUT(C1_DATA4_6) );
  OAI21 U170 ( .IN1(n201), .IN2(n407), .IN3(DP_OP_989_183_2805_n23), .OUT(n106) );
  INVX1 U171 ( .IN(n106), .OUT(C1_DATA11_1) );
  INVX1 U172 ( .IN(DP_OP_981J1_124_6202_n61), .OUT(n107) );
  NAND2X1 U173 ( .IN1(n253), .IN2(DP_OP_981J1_124_6202_n57), .OUT(n108) );
  MUX2X1 U174 ( .IN1(DP_OP_981J1_124_6202_n61), .IN2(n107), .S(n108), .OUT(
        N146) );
  NAND3X1 U175 ( .IN1(n1212), .IN2(n526), .IN3(n927), .OUT(n114) );
  INVX1 U176 ( .IN(n114), .OUT(n115) );
  NAND3X1 U177 ( .IN1(n936), .IN2(n1008), .IN3(n115), .OUT(n1498) );
  INVX1 U178 ( .IN(DP_OP_979_173_2805_n79), .OUT(n125) );
  NOR2X1 U179 ( .IN1(DP_OP_979_173_2805_n1), .IN2(DP_OP_979_173_2805_n39), 
        .OUT(n126) );
  MUX2X1 U180 ( .IN1(DP_OP_979_173_2805_n79), .IN2(n125), .S(n126), .OUT(n127)
         );
  NAND2X1 U181 ( .IN1(n1197), .IN2(n127), .OUT(n1160) );
  NAND2X1 U182 ( .IN1(n417), .IN2(n1378), .OUT(n128) );
  NAND2X1 U183 ( .IN1(n1348), .IN2(n128), .OUT(n1444) );
  NAND3X1 U184 ( .IN1(add_x_35_A_6_), .IN2(n1547), .IN3(add_x_35_A_7_), .OUT(
        n1561) );
  INVX1 U185 ( .IN(DP_OP_981J1_124_6202_n11), .OUT(n129) );
  INVX1 U186 ( .IN(n225), .OUT(n130) );
  AOI22 U187 ( .IN1(n250), .IN2(DP_OP_982J1_125_6202_n175), .IN3(n129), .IN4(
        n130), .OUT(N362) );
  NOR2X1 U188 ( .IN1(n557), .IN2(n639), .OUT(n131) );
  INVX1 U189 ( .IN(n673), .OUT(n132) );
  NAND2X1 U190 ( .IN1(n680), .IN2(n131), .OUT(n133) );
  OAI21 U191 ( .IN1(n367), .IN2(n132), .IN3(n133), .OUT(n867) );
  OAI21 U192 ( .IN1(DP_OP_990_184_2805_n2), .IN2(DP_OP_979_173_2805_n80), 
        .IN3(DP_OP_990_184_2805_n5), .OUT(n134) );
  INVX1 U193 ( .IN(n1272), .OUT(n135) );
  NAND2X1 U194 ( .IN1(DP_OP_989_183_2805_n3), .IN2(DP_OP_989_183_2805_n4), 
        .OUT(n136) );
  NAND2X1 U195 ( .IN1(DP_OP_991_185_2805_n3), .IN2(DP_OP_991_185_2805_n4), 
        .OUT(n137) );
  AOI22 U196 ( .IN1(n1199), .IN2(n136), .IN3(n1198), .IN4(n137), .OUT(n138) );
  OAI21 U197 ( .IN1(n134), .IN2(n135), .IN3(n138), .OUT(n349) );
  AOI22 U198 ( .IN1(n307), .IN2(carry_reg), .IN3(n303), .IN4(n277), .OUT(n139)
         );
  INVX4 U199 ( .IN(n139), .OUT(n538) );
  NOR2X1 U200 ( .IN1(n184), .IN2(n1104), .OUT(n140) );
  INVX1 U201 ( .IN(n140), .OUT(n1097) );
  OAI21 U202 ( .IN1(n284), .IN2(DP_OP_982J1_125_6202_n104), .IN3(n289), .OUT(
        n141) );
  NAND2X1 U203 ( .IN1(DP_OP_982J1_125_6202_n73), .IN2(n141), .OUT(n260) );
  AOI21 U204 ( .IN1(DP_OP_979_173_2805_n78), .IN2(DP_OP_985_179_8739_n30), 
        .IN3(DP_OP_985_179_8739_n11), .OUT(n1122) );
  OAI21 U205 ( .IN1(DP_OP_987_181_8739_n32), .IN2(DP_OP_979_173_2805_n76), 
        .IN3(DP_OP_987_181_8739_n19), .OUT(n142) );
  INVX1 U206 ( .IN(n142), .OUT(C1_DATA9_3) );
  OAI21 U207 ( .IN1(n203), .IN2(n411), .IN3(DP_OP_992_186_8739_n23), .OUT(n143) );
  INVX1 U208 ( .IN(n143), .OUT(C1_DATA7_2) );
  AOI21 U209 ( .IN1(n237), .IN2(n252), .IN3(n247), .OUT(n144) );
  INVX1 U210 ( .IN(n144), .OUT(DP_OP_981J1_124_6202_n106) );
  INVX1 U211 ( .IN(n600), .OUT(n145) );
  NOR2X1 U212 ( .IN1(n380), .IN2(n145), .OUT(n379) );
  AOI21 U213 ( .IN1(DP_OP_979_173_2805_n77), .IN2(DP_OP_979_173_2805_n76), 
        .IN3(DP_OP_986_180_8739_n15), .OUT(n146) );
  INVX1 U214 ( .IN(n146), .OUT(n147) );
  AOI21 U215 ( .IN1(n148), .IN2(n149), .IN3(DP_OP_981_175_8739_n13), .OUT(n150) );
  AOI22 U216 ( .IN1(n1188), .IN2(n147), .IN3(n1187), .IN4(n150), .OUT(n1171)
         );
  INVX1 U217 ( .IN(DP_OP_981_175_8739_n15), .OUT(n148) );
  INVX1 U218 ( .IN(DP_OP_979_173_2805_n77), .OUT(n149) );
  NAND3X1 U219 ( .IN1(DP_OP_982J1_125_6202_n84), .IN2(DP_OP_982J1_125_6202_n83), .IN3(DP_OP_982J1_125_6202_n78), .OUT(n151) );
  NOR2X1 U220 ( .IN1(N422), .IN2(n151), .OUT(n152) );
  NAND2X1 U221 ( .IN1(DP_OP_982J1_125_6202_n77), .IN2(n152), .OUT(n401) );
  NAND3X1 U222 ( .IN1(DP_OP_981J1_124_6202_n77), .IN2(DP_OP_981J1_124_6202_n78), .IN3(n749), .OUT(n153) );
  INVX1 U223 ( .IN(n153), .OUT(n751) );
  INVX1 U224 ( .IN(DP_OP_981J1_124_6202_n99), .OUT(n154) );
  MUX2X1 U225 ( .IN1(n154), .IN2(DP_OP_981J1_124_6202_n99), .S(
        DP_OP_981J1_124_6202_n122), .OUT(N364) );
  AOI21 U226 ( .IN1(DP_OP_979_173_2805_n79), .IN2(DP_OP_984_178_8739_n25), 
        .IN3(DP_OP_984_178_8739_n7), .OUT(n155) );
  INVX1 U227 ( .IN(n155), .OUT(n156) );
  OAI21 U228 ( .IN1(DP_OP_979_173_2805_n79), .IN2(DP_OP_992_186_8739_n29), 
        .IN3(DP_OP_992_186_8739_n7), .OUT(n157) );
  INVX1 U229 ( .IN(n157), .OUT(n158) );
  AOI22 U230 ( .IN1(n1181), .IN2(n156), .IN3(n1271), .IN4(n158), .OUT(n1155)
         );
  AOI21 U231 ( .IN1(DP_OP_979_173_2805_n79), .IN2(DP_OP_986_180_8739_n17), 
        .IN3(DP_OP_986_180_8739_n7), .OUT(n159) );
  INVX1 U232 ( .IN(n159), .OUT(C1_DATA8_6) );
  INVX1 U233 ( .IN(DP_OP_990_184_2805_n51), .OUT(n160) );
  INVX1 U234 ( .IN(DP_OP_979_173_2805_n76), .OUT(n161) );
  AOI22 U235 ( .IN1(DP_OP_979_173_2805_n76), .IN2(n160), .IN3(
        DP_OP_990_184_2805_n51), .IN4(n161), .OUT(C1_DATA12_3) );
  OAI21 U236 ( .IN1(n201), .IN2(n407), .IN3(DP_OP_989_183_2805_n23), .OUT(n162) );
  INVX1 U237 ( .IN(n162), .OUT(C1_DATA13_1) );
  NAND2X1 U238 ( .IN1(n270), .IN2(n267), .OUT(n163) );
  INVX1 U239 ( .IN(n163), .OUT(N420) );
  OAI21 U240 ( .IN1(DP_OP_989_183_2805_n38), .IN2(DP_OP_979_173_2805_n79), 
        .IN3(DP_OP_989_183_2805_n8), .OUT(n164) );
  INVX1 U241 ( .IN(n164), .OUT(n165) );
  INVX1 U242 ( .IN(DP_OP_979_173_2805_n79), .OUT(n166) );
  MUX2X1 U243 ( .IN1(DP_OP_979_173_2805_n79), .IN2(n166), .S(
        DP_OP_991_185_2805_n38), .OUT(n167) );
  AOI22 U244 ( .IN1(n1199), .IN2(n165), .IN3(n1198), .IN4(n167), .OUT(n1163)
         );
  AOI22 U245 ( .IN1(N419), .IN2(Datain1[3]), .IN3(n1411), .IN4(Datain1[1]), 
        .OUT(n168) );
  INVX1 U246 ( .IN(n168), .OUT(n169) );
  NAND2X1 U247 ( .IN1(n1446), .IN2(n169), .OUT(n1371) );
  NAND2X1 U248 ( .IN1(DP_OP_981J1_124_6202_n33), .IN2(DP_OP_981J1_124_6202_n37), .OUT(n170) );
  OAI21 U249 ( .IN1(DP_OP_981J1_124_6202_n33), .IN2(DP_OP_981J1_124_6202_n37), 
        .IN3(n170), .OUT(n325) );
  INVX1 U250 ( .IN(DP_OP_982J1_125_6202_n61), .OUT(n171) );
  NAND2X1 U251 ( .IN1(DP_OP_982J1_125_6202_n56), .IN2(DP_OP_982J1_125_6202_n57), .OUT(n172) );
  MUX2X1 U252 ( .IN1(DP_OP_982J1_125_6202_n61), .IN2(n171), .S(n172), .OUT(
        N158) );
  MUX2X1 U253 ( .IN1(n1293), .IN2(n1292), .S(n1291), .OUT(n173) );
  AOI21 U254 ( .IN1(n1295), .IN2(n1294), .IN3(n173), .OUT(n1302) );
  NOR2X1 U255 ( .IN1(Dataout_valid_BAR), .IN2(n1538), .OUT(n174) );
  INVX1 U256 ( .IN(n174), .OUT(n1539) );
  NOR2X1 U257 ( .IN1(n193), .IN2(n1045), .OUT(n175) );
  INVX1 U258 ( .IN(n175), .OUT(n1096) );
  NOR2X1 U259 ( .IN1(Op2_Mantissa_reg_7_), .IN2(n1561), .OUT(n176) );
  AOI21 U260 ( .IN1(n176), .IN2(n177), .IN3(n178), .OUT(n124) );
  INVX1 U261 ( .IN(n1560), .OUT(n177) );
  INVX1 U262 ( .IN(n1562), .OUT(n178) );
  NAND3X1 U263 ( .IN1(n900), .IN2(n898), .IN3(n899), .OUT(n179) );
  AOI21 U264 ( .IN1(n901), .IN2(n902), .IN3(n179), .OUT(n180) );
  OAI21 U265 ( .IN1(n904), .IN2(n1510), .IN3(n903), .OUT(n181) );
  NAND3X1 U266 ( .IN1(n180), .IN2(n905), .IN3(n181), .OUT(n182) );
  AOI22 U267 ( .IN1(Final_Mantissa_reg[10]), .IN2(n906), .IN3(n429), .IN4(n182), .OUT(n183) );
  INVX1 U268 ( .IN(n183), .OUT(n1062) );
  NAND2X1 U269 ( .IN1(n452), .IN2(n451), .OUT(n453) );
  NANDX2 U270 ( .IN1(n1003), .IN2(n1238), .OUT(n1025) );
  NAND2X1 U271 ( .IN1(n334), .IN2(n487), .OUT(n336) );
  NANDX2 U272 ( .IN1(n962), .IN2(n1500), .OUT(n963) );
  INVX8 U273 ( .IN(Datain2[8]), .OUT(DP_OP_981J1_124_6202_n140) );
  NAND2X1 U274 ( .IN1(n237), .IN2(n245), .OUT(n246) );
  NAND2X1 U275 ( .IN1(n751), .IN2(n750), .OUT(n752) );
  NAND2X1 U276 ( .IN1(n220), .IN2(DP_OP_981J1_124_6202_n140), .OUT(n258) );
  NAND2X1 U277 ( .IN1(DP_OP_981J1_124_6202_n140), .IN2(Datain1[8]), .OUT(
        DP_OP_981J1_124_6202_n124) );
  BUF4X U278 ( .IN(Final_Mantissa_reg[6]), .OUT(n422) );
  NOR2X1 U279 ( .IN1(DP_OP_981J1_124_6202_n20), .IN2(DP_OP_981J1_124_6202_n45), 
        .OUT(n190) );
  NOR2X1 U280 ( .IN1(DP_OP_982J1_125_6202_n20), .IN2(DP_OP_982J1_125_6202_n45), 
        .OUT(n191) );
  NAND2X1 U281 ( .IN1(n1031), .IN2(n1030), .OUT(n1032) );
  INVX4 U282 ( .IN(n1013), .OUT(n981) );
  INVX1 U283 ( .IN(n487), .OUT(n192) );
  NANDX2 U284 ( .IN1(n1046), .IN2(n1047), .OUT(n193) );
  NAND2X1 U285 ( .IN1(n457), .IN2(n456), .OUT(n950) );
  INVX1 U286 ( .IN(DP_OP_982J1_125_6202_n122), .OUT(n269) );
  BUF4X U287 ( .IN(n489), .OUT(n194) );
  NANDX2 U288 ( .IN1(n1143), .IN2(n1142), .OUT(n195) );
  NANDX2 U289 ( .IN1(n196), .IN2(n1141), .OUT(n1144) );
  INVX4 U290 ( .IN(n195), .OUT(n196) );
  INVX4 U291 ( .IN(n1144), .OUT(n1146) );
  INVX1 U292 ( .IN(n410), .OUT(n396) );
  BUF8X U293 ( .IN(Final_Mantissa_reg[1]), .OUT(n427) );
  NAND2X1 U294 ( .IN1(n427), .IN2(n935), .OUT(n1493) );
  BUF8X U295 ( .IN(Final_Mantissa_reg[2]), .OUT(n428) );
  NAND2X1 U296 ( .IN1(n428), .IN2(n535), .OUT(n548) );
  NAND2X1 U297 ( .IN1(n428), .IN2(n477), .OUT(n480) );
  INVX4 U298 ( .IN(n1500), .OUT(n1238) );
  NANDX2 U299 ( .IN1(n1500), .IN2(n965), .OUT(n366) );
  NAND2X1 U300 ( .IN1(n1500), .IN2(n464), .OUT(n465) );
  INVX1 U301 ( .IN(n1530), .OUT(n578) );
  NANDX2 U302 ( .IN1(n1000), .IN2(n1016), .OUT(n1001) );
  NANDX2 U303 ( .IN1(n1272), .IN2(n340), .OUT(n339) );
  INVX4 U304 ( .IN(n1418), .OUT(n1419) );
  INVX8 U305 ( .IN(n1388), .OUT(n197) );
  INVX4 U306 ( .IN(n202), .OUT(n198) );
  NANDX2 U307 ( .IN1(n406), .IN2(n1230), .OUT(n942) );
  NANDX2 U308 ( .IN1(n204), .IN2(DP_OP_982J1_125_6202_n100), .OUT(n271) );
  INVX1 U309 ( .IN(n473), .OUT(n381) );
  NAND2X1 U310 ( .IN1(n500), .IN2(n471), .OUT(n473) );
  NANDX2 U311 ( .IN1(n314), .IN2(n527), .OUT(n928) );
  INVX4 U312 ( .IN(n252), .OUT(n239) );
  INVX4 U313 ( .IN(DP_OP_982J1_125_6202_n66), .OUT(n204) );
  INVX1 U314 ( .IN(n1529), .OUT(Debug[2]) );
  NANDX2 U315 ( .IN1(Datain1[14]), .IN2(n209), .OUT(n436) );
  INVX4 U316 ( .IN(n761), .OUT(n762) );
  INVX1 U317 ( .IN(n418), .OUT(n1314) );
  INVX1 U318 ( .IN(n333), .OUT(n329) );
  NANDX2 U319 ( .IN1(n406), .IN2(n293), .OUT(DP_OP_980_174_8739_n28) );
  NAND2X1 U320 ( .IN1(n312), .IN2(n308), .OUT(n333) );
  INVX4 U321 ( .IN(DP_OP_979_173_2805_n78), .OUT(n199) );
  INVX4 U322 ( .IN(n225), .OUT(n200) );
  NAND2X1 U323 ( .IN1(n868), .IN2(n867), .OUT(n869) );
  NAND2X1 U324 ( .IN1(n602), .IN2(n601), .OUT(n603) );
  NAND2X1 U325 ( .IN1(n675), .IN2(n674), .OUT(n676) );
  NAND2X1 U326 ( .IN1(n573), .IN2(n572), .OUT(n574) );
  NAND2X1 U327 ( .IN1(n625), .IN2(n624), .OUT(n626) );
  INVX1 U328 ( .IN(n1295), .OUT(n1293) );
  NAND2X1 U329 ( .IN1(n1432), .IN2(n1431), .OUT(n1077) );
  INVX1 U330 ( .IN(n1127), .OUT(n1129) );
  INVX1 U331 ( .IN(n1159), .OUT(n1161) );
  INVX1 U332 ( .IN(n1054), .OUT(n1056) );
  NANDX2 U333 ( .IN1(n1510), .IN2(n1484), .OUT(n501) );
  NANDX2 U334 ( .IN1(n1448), .IN2(n1447), .OUT(n1075) );
  NANDX2 U335 ( .IN1(n1337), .IN2(n1336), .OUT(n1338) );
  NAND2X1 U336 ( .IN1(n197), .IN2(n1453), .OUT(n825) );
  NANDX2 U337 ( .IN1(n1370), .IN2(n1446), .OUT(n1412) );
  NAND2X1 U338 ( .IN1(n1197), .IN2(C1_DATA1_3), .OUT(n1055) );
  NANDX2 U339 ( .IN1(n1436), .IN2(n1446), .OUT(n1437) );
  NANDX2 U340 ( .IN1(n1279), .IN2(n1278), .OUT(n1280) );
  INVX1 U341 ( .IN(n1508), .OUT(n1511) );
  NANDX2 U342 ( .IN1(n414), .IN2(n577), .OUT(n1530) );
  INVX1 U343 ( .IN(n1361), .OUT(n1389) );
  NANDX2 U344 ( .IN1(n1249), .IN2(n1248), .OUT(n1250) );
  NAND2X1 U345 ( .IN1(n980), .IN2(n967), .OUT(n968) );
  NAND2X1 U346 ( .IN1(n363), .IN2(n989), .OUT(n990) );
  INVX1 U347 ( .IN(n1026), .OUT(n1015) );
  INVX1 U348 ( .IN(n1399), .OUT(n1400) );
  INVX1 U349 ( .IN(n1329), .OUT(n1335) );
  INVX1 U350 ( .IN(n644), .OUT(n659) );
  NAND2X1 U351 ( .IN1(n681), .IN2(n886), .OUT(n569) );
  NAND2X1 U352 ( .IN1(N419), .IN2(n1406), .OUT(n383) );
  INVX4 U353 ( .IN(n1318), .OUT(n1564) );
  NAND2X1 U354 ( .IN1(n612), .IN2(n611), .OUT(n613) );
  NAND2X1 U355 ( .IN1(n1354), .IN2(n197), .OUT(n1355) );
  NAND2X1 U356 ( .IN1(n1387), .IN2(n356), .OUT(n354) );
  INVX1 U357 ( .IN(n357), .OUT(n356) );
  NAND2X1 U358 ( .IN1(n1498), .IN2(n1482), .OUT(n528) );
  NAND2X1 U359 ( .IN1(DP_OP_982J1_125_6202_n33), .IN2(n255), .OUT(
        DP_OP_982J1_125_6202_n27) );
  INVX4 U360 ( .IN(n395), .OUT(n201) );
  NANDX2 U361 ( .IN1(n1202), .IN2(n1251), .OUT(n1207) );
  INVX1 U362 ( .IN(n919), .OUT(N2921) );
  INVX1 U363 ( .IN(n1493), .OUT(n1204) );
  INVX1 U364 ( .IN(n1008), .OUT(n1201) );
  NANDX2 U365 ( .IN1(DP_OP_981J1_124_6202_n98), .IN2(n235), .OUT(
        DP_OP_981J1_124_6202_n83) );
  NAND2X1 U366 ( .IN1(DP_OP_982J1_125_6202_n33), .IN2(DP_OP_982J1_125_6202_n37), .OUT(n255) );
  NANDX2 U367 ( .IN1(DP_OP_981J1_124_6202_n117), .IN2(n235), .OUT(
        DP_OP_981J1_124_6202_n84) );
  NAND2X1 U368 ( .IN1(n417), .IN2(n198), .OUT(n1349) );
  NANDX2 U369 ( .IN1(n421), .IN2(n694), .OUT(n553) );
  NAND2X1 U370 ( .IN1(n891), .IN2(n583), .OUT(n591) );
  INVX1 U371 ( .IN(n588), .OUT(n589) );
  NANDX2 U372 ( .IN1(n936), .IN2(n518), .OUT(n1519) );
  NANDX2 U373 ( .IN1(n258), .IN2(n256), .OUT(DP_OP_982J1_125_6202_n31) );
  INVX1 U374 ( .IN(n1041), .OUT(n971) );
  NANDX2 U375 ( .IN1(DP_OP_981J1_124_6202_n11), .IN2(n236), .OUT(
        DP_OP_981J1_124_6202_n89) );
  INVX1 U376 ( .IN(n433), .OUT(n1103) );
  INVX1 U377 ( .IN(n893), .OUT(n583) );
  INVX1 U378 ( .IN(n370), .OUT(n372) );
  INVX4 U379 ( .IN(n1203), .OUT(n1229) );
  INVX1 U380 ( .IN(n1489), .OUT(n1490) );
  NANDX2 U381 ( .IN1(n230), .IN2(n228), .OUT(DP_OP_981J1_124_6202_n31) );
  NAND2X1 U382 ( .IN1(n901), .IN2(n1517), .OUT(n875) );
  INVX1 U383 ( .IN(n1387), .OUT(n355) );
  NANDX2 U384 ( .IN1(DP_OP_981J1_124_6202_n11), .IN2(DP_OP_981J1_124_6202_n100), .OUT(n236) );
  NANDX2 U385 ( .IN1(n258), .IN2(DP_OP_982J1_125_6202_n44), .OUT(n256) );
  INVX1 U386 ( .IN(n517), .OUT(n518) );
  INVX1 U387 ( .IN(n1212), .OUT(n941) );
  INVX1 U388 ( .IN(n1584), .OUT(n1296) );
  INVX1 U389 ( .IN(n1578), .OUT(n1579) );
  NAND2X1 U390 ( .IN1(DP_OP_981J1_124_6202_n131), .IN2(n241), .OUT(n242) );
  NAND2X1 U391 ( .IN1(n901), .IN2(n976), .OUT(n539) );
  NANDX2 U392 ( .IN1(n230), .IN2(DP_OP_981J1_124_6202_n44), .OUT(n228) );
  NAND2X1 U393 ( .IN1(n977), .IN2(n976), .OUT(n978) );
  NANDX2 U394 ( .IN1(n1548), .IN2(n1264), .OUT(n1223) );
  INVX1 U395 ( .IN(n1433), .OUT(ExcCheck_Datain_3_) );
  INVX1 U396 ( .IN(n1416), .OUT(ExcCheck_Datain_2_) );
  INVX1 U397 ( .IN(n1374), .OUT(ExcCheck_Datain_1_) );
  INVX1 U398 ( .IN(n1344), .OUT(ExcCheck_Datain_0_) );
  NAND2X1 U399 ( .IN1(n548), .IN2(n1563), .OUT(n549) );
  INVX1 U400 ( .IN(n1440), .OUT(ExcCheck_Datain_4_) );
  NANDX2 U401 ( .IN1(n1556), .IN2(n1264), .OUT(n1274) );
  INVX1 U402 ( .IN(n1461), .OUT(ExcCheck_Datain_6_) );
  INVX1 U403 ( .IN(n1449), .OUT(ExcCheck_Datain_5_) );
  NANDX2 U404 ( .IN1(n422), .IN2(n1520), .OUT(n1492) );
  INVX1 U405 ( .IN(n253), .OUT(DP_OP_982J1_125_6202_n16) );
  NAND2X1 U406 ( .IN1(DP_OP_981J1_124_6202_n127), .IN2(n237), .OUT(n248) );
  INVX1 U407 ( .IN(DP_OP_981J1_124_6202_n124), .OUT(n243) );
  INVX1 U408 ( .IN(n906), .OUT(n911) );
  NAND2X1 U409 ( .IN1(n1556), .IN2(n506), .OUT(n508) );
  INVX4 U410 ( .IN(n506), .OUT(n1264) );
  INVX1 U411 ( .IN(DP_OP_982J1_125_6202_n56), .OUT(DP_OP_981J1_124_6202_n16)
         );
  NAND2X1 U412 ( .IN1(n429), .IN2(n436), .OUT(n437) );
  NAND2X1 U413 ( .IN1(n697), .IN2(n431), .OUT(n909) );
  NANDX2 U414 ( .IN1(n1309), .IN2(n1308), .OUT(n1535) );
  INVX1 U415 ( .IN(DP_OP_981J1_124_6202_n121), .OUT(DP_OP_981J1_124_6202_n119)
         );
  INVX1 U416 ( .IN(n1589), .OUT(Debug[4]) );
  INVX1 U417 ( .IN(n1516), .OUT(Debug[1]) );
  INVX1 U418 ( .IN(n1486), .OUT(Debug[0]) );
  INVX4 U419 ( .IN(DP_OP_985_179_8739_n27), .OUT(n203) );
  NANDX2 U420 ( .IN1(n425), .IN2(n1488), .OUT(n927) );
  NAND2X1 U421 ( .IN1(n1626), .IN2(n429), .OUT(n1628) );
  INVX1 U422 ( .IN(n1626), .OUT(n431) );
  NANDX2 U423 ( .IN1(StateMC[2]), .IN2(n1305), .OUT(Dataout_valid_BAR) );
  NANDX2 U424 ( .IN1(Datain1[10]), .IN2(n1570), .OUT(DP_OP_982J1_125_6202_n130) );
  NAND2X1 U425 ( .IN1(n186), .IN2(n297), .OUT(n448) );
  INVX4 U426 ( .IN(n1556), .OUT(n1548) );
  INVX1 U427 ( .IN(DP_OP_982J1_125_6202_n112), .OUT(DP_OP_982J1_125_6202_n129)
         );
  INVX1 U428 ( .IN(n1619), .OUT(n1331) );
  INVX4 U429 ( .IN(DP_OP_987_181_8739_n27), .OUT(n205) );
  NANDX2 U430 ( .IN1(n429), .IN2(n1563), .OUT(n1308) );
  NAND2X1 U431 ( .IN1(n429), .IN2(n550), .OUT(n1309) );
  NANDX2 U432 ( .IN1(n424), .IN2(n296), .OUT(n1219) );
  INVX1 U433 ( .IN(DP_OP_982J1_125_6202_n181), .OUT(DP_OP_981J1_124_6202_n135)
         );
  NAND2X1 U434 ( .IN1(n419), .IN2(n420), .OUT(n536) );
  INVX1 U435 ( .IN(n416), .OUT(n1376) );
  NANDX2 U436 ( .IN1(n300), .IN2(n1566), .OUT(n1581) );
  NANDX2 U437 ( .IN1(Debug_reg[3]), .IN2(n1588), .OUT(n1537) );
  INVX4 U438 ( .IN(DP_OP_982J1_125_6202_n180), .OUT(n206) );
  INVX4 U439 ( .IN(DP_OP_979_173_2805_n77), .OUT(n207) );
  INVX4 U440 ( .IN(DP_OP_982J1_125_6202_n182), .OUT(n209) );
  INVX4 U441 ( .IN(DP_OP_980_174_8739_n28), .OUT(n210) );
  BUF4X U442 ( .IN(Datain1[7]), .OUT(n225) );
  NAND2X1 U443 ( .IN1(n296), .IN2(n310), .OUT(n509) );
  NANDX2 U444 ( .IN1(add_x_35_A_0_), .IN2(add_x_35_A_1_), .OUT(n1479) );
  INVX8 U445 ( .IN(DP_OP_982J1_125_6202_n177), .OUT(n220) );
  BUF4X U446 ( .IN(Final_Mantissa_reg[7]), .OUT(n423) );
  NANDX2 U447 ( .IN1(n1003), .IN2(n1002), .OUT(n1004) );
  INVX1 U448 ( .IN(n963), .OUT(n964) );
  INVX1 U449 ( .IN(n1110), .OUT(n1112) );
  INVX1 U450 ( .IN(n1022), .OUT(n1034) );
  MUX2X1 U451 ( .IN1(n424), .IN2(n310), .S(n488), .OUT(n221) );
  MUX2X1 U452 ( .IN1(n310), .IN2(n424), .S(n488), .OUT(n224) );
  INVX1 U453 ( .IN(n495), .OUT(n496) );
  NAND2X1 U454 ( .IN1(DP_OP_979_173_2805_n48), .IN2(DP_OP_979_173_2805_n77), 
        .OUT(DP_OP_979_173_2805_n14) );
  INVX4 U455 ( .IN(n204), .OUT(n226) );
  BUF4X U456 ( .IN(N362), .OUT(N147) );
  AOI21 U457 ( .IN1(DP_OP_981J1_124_6202_n131), .IN2(n243), .IN3(
        DP_OP_981J1_124_6202_n119), .OUT(n244) );
  OAI21 U458 ( .IN1(DP_OP_981J1_124_6202_n117), .IN2(DP_OP_981J1_124_6202_n17), 
        .IN3(DP_OP_982J1_125_6202_n130), .OUT(DP_OP_981J1_124_6202_n114) );
  OAI21 U459 ( .IN1(DP_OP_981J1_124_6202_n123), .IN2(DP_OP_981J1_124_6202_n11), 
        .IN3(DP_OP_981J1_124_6202_n124), .OUT(DP_OP_981J1_124_6202_n122) );
  OAI21 U460 ( .IN1(DP_OP_981J1_124_6202_n11), .IN2(n242), .IN3(n244), .OUT(
        n245) );
  OAI21 U461 ( .IN1(n238), .IN2(DP_OP_981J1_124_6202_n117), .IN3(n239), .OUT(
        n240) );
  OAI21 U462 ( .IN1(n248), .IN2(n239), .IN3(DP_OP_981J1_124_6202_n105), .OUT(
        n249) );
  AOI21 U463 ( .IN1(n247), .IN2(DP_OP_981J1_124_6202_n127), .IN3(n249), .OUT(
        DP_OP_981J1_124_6202_n101) );
  OAI21 U464 ( .IN1(n238), .IN2(n246), .IN3(DP_OP_981J1_124_6202_n108), .OUT(
        n247) );
  INVX4 U465 ( .IN(n250), .OUT(DP_OP_981J1_124_6202_n11) );
  OAI21 U466 ( .IN1(n234), .IN2(n233), .IN3(n251), .OUT(N366) );
  OAI21 U467 ( .IN1(DP_OP_981J1_124_6202_n112), .IN2(DP_OP_982J1_125_6202_n130), .IN3(DP_OP_981J1_124_6202_n113), .OUT(n252) );
  INVX1 U468 ( .IN(DP_OP_981J1_124_6202_n123), .OUT(n241) );
  INVX1 U469 ( .IN(Datain2[11]), .OUT(DP_OP_981J1_124_6202_n137) );
  INVX1 U470 ( .IN(DP_OP_981J1_124_6202_n112), .OUT(DP_OP_981J1_124_6202_n129)
         );
  INVX1 U471 ( .IN(DP_OP_981J1_124_6202_n101), .OUT(n231) );
  NAND2X1 U472 ( .IN1(n272), .IN2(n230), .OUT(n229) );
  INVX1 U473 ( .IN(n229), .OUT(DP_OP_981J1_124_6202_n45) );
  NAND2X1 U474 ( .IN1(DP_OP_981J1_124_6202_n44), .IN2(n228), .OUT(
        DP_OP_981J1_124_6202_n4) );
  NAND2X1 U475 ( .IN1(n1570), .IN2(DP_OP_982J1_125_6202_n130), .OUT(
        DP_OP_981J1_124_6202_n57) );
  NANDX2 U476 ( .IN1(DP_OP_982J1_125_6202_n175), .IN2(n200), .OUT(n250) );
  INVX4 U477 ( .IN(DP_OP_981J1_124_6202_n120), .OUT(DP_OP_981J1_124_6202_n131)
         );
  INVX4 U478 ( .IN(n245), .OUT(DP_OP_981J1_124_6202_n117) );
  INVX4 U479 ( .IN(DP_OP_982J1_125_6202_n58), .OUT(DP_OP_981J1_124_6202_n17)
         );
  INVX4 U480 ( .IN(DP_OP_981J1_124_6202_n114), .OUT(n234) );
  INVX4 U481 ( .IN(DP_OP_981J1_124_6202_n97), .OUT(n233) );
  NANDX2 U482 ( .IN1(n233), .IN2(n234), .OUT(n251) );
  NANDX2 U483 ( .IN1(DP_OP_981J1_124_6202_n98), .IN2(DP_OP_981J1_124_6202_n117), .OUT(n235) );
  INVX4 U484 ( .IN(n240), .OUT(DP_OP_981J1_124_6202_n109) );
  INVX4 U485 ( .IN(DP_OP_981J1_124_6202_n107), .OUT(n237) );
  NANDX2 U486 ( .IN1(DP_OP_981J1_124_6202_n96), .IN2(DP_OP_981J1_124_6202_n109), .OUT(n232) );
  NANDX2 U487 ( .IN1(DP_OP_981J1_124_6202_n109), .IN2(n232), .OUT(
        DP_OP_981J1_124_6202_n78) );
  INVX4 U488 ( .IN(DP_OP_981J1_124_6202_n104), .OUT(DP_OP_981J1_124_6202_n127)
         );
  NANDX2 U489 ( .IN1(DP_OP_982J1_125_6202_n139), .IN2(n272), .OUT(n230) );
  INVX4 U490 ( .IN(n227), .OUT(DP_OP_981J1_124_6202_n20) );
  INVX4 U491 ( .IN(DP_OP_981J1_124_6202_n8), .OUT(N151) );
  NANDX2 U492 ( .IN1(DP_OP_981J1_124_6202_n96), .IN2(n232), .OUT(
        DP_OP_981J1_124_6202_n77) );
  NANDX2 U493 ( .IN1(DP_OP_982J1_125_6202_n139), .IN2(n230), .OUT(n227) );
  NAND2X1 U494 ( .IN1(DP_OP_981J1_124_6202_n100), .IN2(n236), .OUT(
        DP_OP_981J1_124_6202_n90) );
  INVX4 U495 ( .IN(DP_OP_982J1_125_6202_n57), .OUT(DP_OP_981J1_124_6202_n15)
         );
  NANDX2 U496 ( .IN1(DP_OP_981J1_124_6202_n129), .IN2(DP_OP_982J1_125_6202_n58), .OUT(n238) );
  NOR2X1 U497 ( .IN1(DP_OP_982J1_125_6202_n175), .IN2(n204), .OUT(
        DP_OP_982J1_125_6202_n34) );
  NOR2X1 U498 ( .IN1(n200), .IN2(n204), .OUT(DP_OP_982J1_125_6202_n35) );
  INVX1 U499 ( .IN(DP_OP_982J1_125_6202_n123), .OUT(DP_OP_982J1_125_6202_n132)
         );
  NAND2X1 U500 ( .IN1(DP_OP_981J1_124_6202_n140), .IN2(n258), .OUT(n257) );
  INVX1 U501 ( .IN(n257), .OUT(DP_OP_982J1_125_6202_n45) );
  NAND2X1 U502 ( .IN1(n204), .IN2(n271), .OUT(DP_OP_982J1_125_6202_n89) );
  OAI21 U503 ( .IN1(DP_OP_982J1_125_6202_n112), .IN2(DP_OP_982J1_125_6202_n58), 
        .IN3(DP_OP_982J1_125_6202_n113), .OUT(n275) );
  NAND3X1 U504 ( .IN1(DP_OP_982J1_125_6202_n131), .IN2(
        DP_OP_982J1_125_6202_n129), .IN3(DP_OP_982J1_125_6202_n122), .OUT(n280) );
  AOI21 U505 ( .IN1(DP_OP_982J1_125_6202_n122), .IN2(DP_OP_982J1_125_6202_n131), .IN3(DP_OP_982J1_125_6202_n119), .OUT(DP_OP_982J1_125_6202_n117) );
  NANDX2 U506 ( .IN1(n225), .IN2(n281), .OUT(DP_OP_982J1_125_6202_n66) );
  NOR2X1 U507 ( .IN1(n285), .IN2(DP_OP_982J1_125_6202_n128), .OUT(n286) );
  NOR2X1 U508 ( .IN1(n285), .IN2(n283), .OUT(n287) );
  AOI22 U509 ( .IN1(n286), .IN2(n282), .IN3(n287), .IN4(n288), .OUT(n263) );
  OAI21 U510 ( .IN1(DP_OP_982J1_125_6202_n104), .IN2(n284), .IN3(n289), .OUT(
        n261) );
  AOI21 U511 ( .IN1(n284), .IN2(n283), .IN3(DP_OP_982J1_125_6202_n95), .OUT(
        DP_OP_982J1_125_6202_n74) );
  NAND3X1 U512 ( .IN1(DP_OP_982J1_125_6202_n96), .IN2(n291), .IN3(n290), .OUT(
        n264) );
  INVX4 U513 ( .IN(Datain1[8]), .OUT(n272) );
  INVX1 U514 ( .IN(Datain1[11]), .OUT(DP_OP_982J1_125_6202_n137) );
  INVX1 U515 ( .IN(Datain1[10]), .OUT(n259) );
  INVX1 U516 ( .IN(Datain1[12]), .OUT(DP_OP_982J1_125_6202_n136) );
  INVX1 U517 ( .IN(DP_OP_982J1_125_6202_n130), .OUT(n273) );
  NAND2X1 U518 ( .IN1(DP_OP_982J1_125_6202_n117), .IN2(n265), .OUT(
        DP_OP_982J1_125_6202_n84) );
  INVX1 U519 ( .IN(Datain1[13]), .OUT(DP_OP_982J1_125_6202_n135) );
  INVX1 U520 ( .IN(n263), .OUT(DP_OP_982J1_125_6202_n75) );
  NAND2X1 U521 ( .IN1(Datain1[10]), .IN2(DP_OP_982J1_125_6202_n130), .OUT(n253) );
  NAND2X1 U522 ( .IN1(DP_OP_982J1_125_6202_n44), .IN2(n256), .OUT(
        DP_OP_982J1_125_6202_n4) );
  NAND2X1 U523 ( .IN1(n259), .IN2(DP_OP_982J1_125_6202_n58), .OUT(
        DP_OP_982J1_125_6202_n57) );
  NAND2X1 U524 ( .IN1(Datain2[10]), .IN2(DP_OP_982J1_125_6202_n58), .OUT(
        DP_OP_982J1_125_6202_n56) );
  NAND2X1 U525 ( .IN1(DP_OP_982J1_125_6202_n37), .IN2(n255), .OUT(
        DP_OP_982J1_125_6202_n28) );
  INVX4 U526 ( .IN(DP_OP_982J1_125_6202_n175), .OUT(n281) );
  NANDX2 U527 ( .IN1(DP_OP_982J1_125_6202_n100), .IN2(n271), .OUT(
        DP_OP_982J1_125_6202_n90) );
  INVX4 U528 ( .IN(DP_OP_982J1_125_6202_n120), .OUT(DP_OP_982J1_125_6202_n131)
         );
  INVX4 U529 ( .IN(DP_OP_982J1_125_6202_n99), .OUT(n266) );
  NANDX2 U530 ( .IN1(n269), .IN2(n266), .OUT(n268) );
  NANDX2 U531 ( .IN1(n279), .IN2(n280), .OUT(n276) );
  NANDX2 U532 ( .IN1(Datain2[10]), .IN2(n259), .OUT(DP_OP_982J1_125_6202_n58)
         );
  INVX4 U533 ( .IN(n275), .OUT(n291) );
  NANDX2 U534 ( .IN1(n290), .IN2(n291), .OUT(n278) );
  INVX4 U535 ( .IN(n278), .OUT(n288) );
  INVX4 U536 ( .IN(DP_OP_982J1_125_6202_n107), .OUT(DP_OP_982J1_125_6202_n128)
         );
  NANDX2 U537 ( .IN1(DP_OP_982J1_125_6202_n96), .IN2(n264), .OUT(
        DP_OP_982J1_125_6202_n77) );
  NANDX2 U538 ( .IN1(DP_OP_982J1_125_6202_n98), .IN2(DP_OP_982J1_125_6202_n117), .OUT(n265) );
  INVX4 U539 ( .IN(DP_OP_982J1_125_6202_n104), .OUT(DP_OP_982J1_125_6202_n127)
         );
  INVX4 U540 ( .IN(DP_OP_982J1_125_6202_n95), .OUT(n262) );
  INVX4 U541 ( .IN(n282), .OUT(n283) );
  NANDX2 U542 ( .IN1(DP_OP_982J1_125_6202_n128), .IN2(n278), .OUT(n284) );
  NANDX2 U543 ( .IN1(DP_OP_982J1_125_6202_n68), .IN2(DP_OP_982J1_125_6202_n67), 
        .OUT(N425) );
  INVX4 U544 ( .IN(n254), .OUT(DP_OP_982J1_125_6202_n20) );
  INVX4 U545 ( .IN(DP_OP_982J1_125_6202_n12), .OUT(DP_OP_982J1_125_6202_n63)
         );
  INVX4 U546 ( .IN(DP_OP_982J1_125_6202_n8), .OUT(N155) );
  NANDX2 U547 ( .IN1(n269), .IN2(n268), .OUT(n270) );
  NANDX2 U548 ( .IN1(n266), .IN2(n268), .OUT(n267) );
  NANDX2 U549 ( .IN1(n288), .IN2(n264), .OUT(DP_OP_982J1_125_6202_n78) );
  NANDX2 U550 ( .IN1(DP_OP_982J1_125_6202_n108), .IN2(n262), .OUT(n282) );
  NANDX2 U551 ( .IN1(n261), .IN2(n260), .OUT(DP_OP_982J1_125_6202_n68) );
  NANDX2 U552 ( .IN1(DP_OP_982J1_125_6202_n130), .IN2(n276), .OUT(n290) );
  NANDX2 U553 ( .IN1(n220), .IN2(n258), .OUT(n254) );
  INVX4 U554 ( .IN(DP_OP_982J1_125_6202_n108), .OUT(n285) );
  NANDX2 U555 ( .IN1(DP_OP_982J1_125_6202_n73), .IN2(n260), .OUT(
        DP_OP_982J1_125_6202_n67) );
  INVX4 U556 ( .IN(DP_OP_982J1_125_6202_n121), .OUT(DP_OP_982J1_125_6202_n119)
         );
  NANDX2 U557 ( .IN1(DP_OP_982J1_125_6202_n119), .IN2(
        DP_OP_982J1_125_6202_n129), .OUT(n279) );
  INVX4 U558 ( .IN(Datain1[9]), .OUT(DP_OP_982J1_125_6202_n139) );
  NANDX2 U559 ( .IN1(DP_OP_982J1_125_6202_n98), .IN2(n265), .OUT(
        DP_OP_982J1_125_6202_n83) );
  INVX4 U560 ( .IN(DP_OP_981J1_124_6202_n57), .OUT(DP_OP_982J1_125_6202_n15)
         );
  NANDX2 U561 ( .IN1(n883), .IN2(n882), .OUT(n113) );
  NANDX2 U562 ( .IN1(n426), .IN2(n881), .OUT(n882) );
  INVX1 U563 ( .IN(n567), .OUT(n568) );
  NAND2X1 U564 ( .IN1(n426), .IN2(n485), .OUT(n367) );
  NANDX2 U565 ( .IN1(n999), .IN2(n998), .OUT(n1016) );
  NANDX2 U566 ( .IN1(n979), .IN2(n999), .OUT(n983) );
  NAND2X1 U567 ( .IN1(n308), .IN2(n298), .OUT(n447) );
  NANDX2 U568 ( .IN1(n1521), .IN2(n948), .OUT(n999) );
  NANDX2 U569 ( .IN1(DP_OP_979_173_2805_n76), .IN2(Final_Exponent_reg[0]), 
        .OUT(n932) );
  BUF4X U570 ( .IN(N691), .OUT(n426) );
  NAND2X1 U571 ( .IN1(n1373), .IN2(n1372), .OUT(n1079) );
  INVX4 U572 ( .IN(n1369), .OUT(n1379) );
  INVX4 U573 ( .IN(n640), .OUT(n666) );
  NANDX2 U574 ( .IN1(n901), .IN2(n578), .OUT(n640) );
  NANDX2 U575 ( .IN1(n961), .IN2(n960), .OUT(n962) );
  INVX1 U576 ( .IN(n447), .OUT(n443) );
  BUF4X U577 ( .IN(Final_Mantissa_reg[5]), .OUT(n421) );
  INVX1 U578 ( .IN(n526), .OUT(n527) );
  NAND2X1 U579 ( .IN1(n423), .IN2(n1488), .OUT(n526) );
  INVX1 U580 ( .IN(n1304), .OUT(n1305) );
  INVX4 U581 ( .IN(n1499), .OUT(n1532) );
  INVX4 U582 ( .IN(n641), .OUT(n663) );
  INVX4 U583 ( .IN(n500), .OUT(n951) );
  INVX4 U584 ( .IN(n1011), .OUT(n1503) );
  NANDX2 U585 ( .IN1(n314), .IN2(n487), .OUT(n488) );
  NANDX2 U586 ( .IN1(n1003), .IN2(n942), .OUT(n1235) );
  INVX4 U587 ( .IN(RSTn_BAR), .OUT(n429) );
  NANDX2 U588 ( .IN1(n1513), .IN2(n1512), .OUT(n1514) );
  NAND2X1 U589 ( .IN1(n421), .IN2(n537), .OUT(n558) );
  NANDX2 U590 ( .IN1(n1563), .IN2(n908), .OUT(n893) );
  INVX1 U591 ( .IN(n520), .OUT(n524) );
  NANDX2 U592 ( .IN1(n944), .IN2(n352), .OUT(n351) );
  NAND2X1 U593 ( .IN1(n426), .IN2(n299), .OUT(n520) );
  INVX1 U594 ( .IN(n1358), .OUT(n1359) );
  NANDX2 U595 ( .IN1(N362), .IN2(n197), .OUT(n748) );
  NANDX2 U596 ( .IN1(n353), .IN2(n197), .OUT(n1398) );
  INVX4 U597 ( .IN(n354), .OUT(n353) );
  BUF4X U598 ( .IN(n1622), .OUT(n413) );
  INVX1 U599 ( .IN(Datain1[14]), .OUT(n1615) );
  NAND2X1 U600 ( .IN1(n422), .IN2(n559), .OUT(n582) );
  NANDX2 U601 ( .IN1(DP_OP_979_173_2805_n52), .IN2(n201), .OUT(
        DP_OP_989_183_2805_n1) );
  NANDX2 U602 ( .IN1(n965), .IN2(n964), .OUT(n980) );
  NANDX2 U603 ( .IN1(n453), .IN2(n381), .OUT(n380) );
  BUF4X U604 ( .IN(n1509), .OUT(n414) );
  INVX4 U605 ( .IN(n997), .OUT(n944) );
  NAND2X1 U606 ( .IN1(n186), .IN2(n311), .OUT(n515) );
  INVX4 U607 ( .IN(n1350), .OUT(n1377) );
  NANDX2 U608 ( .IN1(N160), .IN2(n775), .OUT(n786) );
  NANDX2 U609 ( .IN1(N148), .IN2(n763), .OUT(n770) );
  NANDX2 U610 ( .IN1(N144), .IN2(n826), .OUT(n839) );
  NANDX2 U611 ( .IN1(N156), .IN2(n803), .OUT(n814) );
  NANDX2 U612 ( .IN1(N152), .IN2(n729), .OUT(n740) );
  NANDX2 U613 ( .IN1(N164), .IN2(n703), .OUT(n714) );
  NANDX2 U614 ( .IN1(n1352), .IN2(n769), .OUT(n1454) );
  INVX1 U615 ( .IN(DP_OP_984_178_8739_n26), .OUT(DP_OP_984_178_8739_n15) );
  INVX4 U616 ( .IN(n693), .OUT(n597) );
  NANDX2 U617 ( .IN1(n1237), .IN2(n1241), .OUT(n921) );
  INVX4 U618 ( .IN(n920), .OUT(n1241) );
  NANDX2 U619 ( .IN1(n194), .IN2(n221), .OUT(n920) );
  NANDX2 U620 ( .IN1(n414), .IN2(n980), .OUT(n1013) );
  NAND2X1 U621 ( .IN1(n423), .IN2(n422), .OUT(n371) );
  NAND2X1 U622 ( .IN1(n423), .IN2(n457), .OUT(n373) );
  NANDX2 U623 ( .IN1(n296), .IN2(n451), .OUT(n489) );
  NANDX2 U624 ( .IN1(Final_Mantissa_reg[10]), .IN2(n450), .OUT(n335) );
  NANDX2 U625 ( .IN1(n1408), .IN2(n1407), .OUT(n1410) );
  INVX4 U626 ( .IN(Datain2[10]), .OUT(n1570) );
  NANDX2 U627 ( .IN1(n436), .IN2(n392), .OUT(n391) );
  BUF4X U628 ( .IN(Datain2[14]), .OUT(DP_OP_982J1_125_6202_n182) );
  NAND2X1 U629 ( .IN1(add_x_35_A_8_), .IN2(add_x_35_A_9_), .OUT(n1560) );
  INVX1 U630 ( .IN(n1441), .OUT(n1442) );
  INVX1 U631 ( .IN(n682), .OUT(n691) );
  NANDX2 U632 ( .IN1(n800), .IN2(n799), .OUT(n403) );
  NANDX2 U633 ( .IN1(n429), .IN2(n1303), .OUT(n922) );
  NAND2X1 U634 ( .IN1(Final_Mantissa_reg[10]), .IN2(n424), .OUT(n892) );
  INVX4 U635 ( .IN(n1220), .OUT(n1221) );
  INVX4 U636 ( .IN(n1200), .OUT(n350) );
  NANDX2 U637 ( .IN1(n1197), .IN2(C1_DATA1_4), .OUT(n1173) );
  NANDX2 U638 ( .IN1(n884), .IN2(n855), .OUT(n874) );
  NANDX2 U639 ( .IN1(n901), .IN2(n1522), .OUT(n484) );
  INVX4 U640 ( .IN(n461), .OUT(n469) );
  INVX4 U641 ( .IN(n497), .OUT(n498) );
  NANDX2 U642 ( .IN1(n1226), .IN2(n496), .OUT(n497) );
  NANDX2 U643 ( .IN1(n1482), .IN2(n530), .OUT(n648) );
  NANDX2 U644 ( .IN1(n1498), .IN2(n531), .OUT(n529) );
  INVX4 U645 ( .IN(n1274), .OUT(n1517) );
  INVX1 U646 ( .IN(DP_OP_988_182_8739_n25), .OUT(DP_OP_988_182_8739_n11) );
  INVX1 U647 ( .IN(DP_OP_987_181_8739_n29), .OUT(DP_OP_987_181_8739_n11) );
  INVX1 U648 ( .IN(DP_OP_981_175_8739_n29), .OUT(DP_OP_981_175_8739_n11) );
  NANDX2 U649 ( .IN1(DP_OP_979_173_2805_n52), .IN2(DP_OP_979_173_2805_n58), 
        .OUT(DP_OP_979_173_2805_n1) );
  NAND2X1 U650 ( .IN1(n1025), .IN2(n1023), .OUT(n1029) );
  NANDX2 U651 ( .IN1(n1227), .IN2(n1278), .OUT(n1010) );
  INVX4 U652 ( .IN(n470), .OUT(n476) );
  NANDX2 U653 ( .IN1(n409), .IN2(DP_OP_981_175_8739_n23), .OUT(
        DP_OP_981_175_8739_n31) );
  NANDX2 U654 ( .IN1(n409), .IN2(DP_OP_984_178_8739_n23), .OUT(
        DP_OP_984_178_8739_n27) );
  NANDX2 U655 ( .IN1(n409), .IN2(DP_OP_992_186_8739_n23), .OUT(
        DP_OP_985_179_8739_n31) );
  INVX4 U656 ( .IN(n465), .OUT(n468) );
  INVX4 U657 ( .IN(n335), .OUT(n334) );
  NAND2X1 U658 ( .IN1(n950), .IN2(n686), .OUT(n952) );
  NANDX2 U659 ( .IN1(n477), .IN2(n332), .OUT(n331) );
  NANDX2 U660 ( .IN1(n362), .IN2(n361), .OUT(n360) );
  INVX4 U661 ( .IN(n427), .OUT(n361) );
  INVX4 U662 ( .IN(n428), .OUT(n362) );
  NANDX2 U663 ( .IN1(n939), .IN2(n938), .OUT(n940) );
  NANDX2 U664 ( .IN1(n1202), .IN2(n975), .OUT(n938) );
  INVX4 U665 ( .IN(n936), .OUT(n1202) );
  INVX1 U666 ( .IN(n933), .OUT(n934) );
  INVX4 U667 ( .IN(n1003), .OUT(n1239) );
  NANDX2 U668 ( .IN1(n293), .IN2(n1230), .OUT(n1003) );
  NANDX2 U669 ( .IN1(n292), .IN2(n1215), .OUT(n1237) );
  INVX4 U670 ( .IN(n1244), .OUT(n1215) );
  NANDX2 U671 ( .IN1(n294), .IN2(n930), .OUT(n992) );
  NANDX2 U672 ( .IN1(n202), .IN2(n1411), .OUT(n1323) );
  INVX4 U673 ( .IN(n383), .OUT(n382) );
  NANDX2 U674 ( .IN1(n1317), .IN2(n1405), .OUT(n1408) );
  NANDX2 U675 ( .IN1(n1319), .IN2(n1405), .OUT(n1320) );
  NANDX2 U676 ( .IN1(n392), .IN2(n389), .OUT(n388) );
  NANDX2 U677 ( .IN1(n418), .IN2(n1378), .OUT(n1450) );
  INVX4 U678 ( .IN(n391), .OUT(n390) );
  INVX4 U679 ( .IN(n1537), .OUT(Debug[3]) );
  NAND2X1 U680 ( .IN1(StateMC[0]), .IN2(StateMC[1]), .OUT(n1304) );
  INVX4 U681 ( .IN(n1474), .OUT(ExcCheck_Datain_14_) );
  INVX4 U682 ( .IN(n1473), .OUT(ExcCheck_Datain_12_) );
  INVX4 U683 ( .IN(n1472), .OUT(ExcCheck_Datain_11_) );
  INVX4 U684 ( .IN(n1470), .OUT(ExcCheck_Datain_9_) );
  INVX4 U685 ( .IN(n1469), .OUT(ExcCheck_Datain_8_) );
  INVX1 U686 ( .IN(Datain2[15]), .OUT(n440) );
  INVX1 U687 ( .IN(Datain1[15]), .OUT(n442) );
  INVX4 U688 ( .IN(n1262), .OUT(n1285) );
  NAND2X1 U689 ( .IN1(Datain1[13]), .IN2(n197), .OUT(n1164) );
  INVX4 U690 ( .IN(n630), .OUT(n634) );
  INVX4 U691 ( .IN(n629), .OUT(n637) );
  NANDX2 U692 ( .IN1(n1435), .IN2(n1451), .OUT(n1438) );
  NANDX2 U693 ( .IN1(n1457), .IN2(n1456), .OUT(n1458) );
  INVX4 U694 ( .IN(n1450), .OUT(n1452) );
  INVX4 U695 ( .IN(n864), .OUT(n1531) );
  INVX4 U696 ( .IN(n1453), .OUT(n1463) );
  NANDX2 U697 ( .IN1(n609), .IN2(n608), .OUT(n630) );
  NANDX2 U698 ( .IN1(n607), .IN2(n606), .OUT(n629) );
  INVX4 U699 ( .IN(n890), .OUT(n552) );
  INVX4 U700 ( .IN(n658), .OUT(n681) );
  INVX4 U701 ( .IN(n905), .OUT(n679) );
  INVX4 U702 ( .IN(n403), .OUT(n402) );
  INVX4 U703 ( .IN(n777), .OUT(n784) );
  INVX4 U704 ( .IN(n774), .OUT(n788) );
  NANDX2 U705 ( .IN1(n773), .IN2(N161), .OUT(n774) );
  INVX4 U706 ( .IN(n765), .OUT(n767) );
  NANDX2 U707 ( .IN1(n1289), .IN2(n1288), .OUT(n1538) );
  NANDX2 U708 ( .IN1(n908), .IN2(n907), .OUT(n1300) );
  INVX4 U709 ( .IN(n1292), .OUT(n1294) );
  NANDX2 U710 ( .IN1(n1254), .IN2(n1253), .OUT(n1284) );
  NANDX2 U711 ( .IN1(n1222), .IN2(n1221), .OUT(n1276) );
  NANDX2 U712 ( .IN1(n1209), .IN2(n1208), .OUT(n1266) );
  INVX4 U713 ( .IN(n1277), .OUT(n1208) );
  NANDX2 U714 ( .IN1(n1207), .IN2(n1206), .OUT(n1277) );
  NANDX2 U715 ( .IN1(n350), .IN2(n347), .OUT(n346) );
  NANDX2 U716 ( .IN1(n295), .IN2(DP_OP_983_177_8739_n11), .OUT(
        DP_OP_983_177_8739_n28) );
  NANDX2 U717 ( .IN1(n1325), .IN2(n1324), .OUT(n1435) );
  NANDX2 U718 ( .IN1(n1315), .IN2(n1325), .OUT(n1436) );
  NANDX2 U719 ( .IN1(n416), .IN2(n1378), .OUT(n1325) );
  NANDX2 U720 ( .IN1(n1314), .IN2(n198), .OUT(n1457) );
  NANDX2 U721 ( .IN1(n337), .IN2(n344), .OUT(n343) );
  INVX4 U722 ( .IN(n338), .OUT(n337) );
  NANDX2 U723 ( .IN1(n1173), .IN2(n1174), .OUT(n338) );
  NAND2X1 U724 ( .IN1(Datain1[11]), .IN2(n197), .OUT(n1177) );
  INVX4 U725 ( .IN(n829), .OUT(n837) );
  INVX4 U726 ( .IN(n805), .OUT(n812) );
  INVX4 U727 ( .IN(n586), .OUT(n688) );
  NANDX2 U728 ( .IN1(n585), .IN2(n584), .OUT(n586) );
  NANDX2 U729 ( .IN1(n580), .IN2(n581), .OUT(n693) );
  INVX4 U730 ( .IN(n731), .OUT(n738) );
  INVX4 U731 ( .IN(n728), .OUT(n742) );
  NANDX2 U732 ( .IN1(n727), .IN2(N153), .OUT(n728) );
  INVX4 U733 ( .IN(n705), .OUT(n712) );
  INVX4 U734 ( .IN(n697), .OUT(n1569) );
  INVX4 U735 ( .IN(n1297), .OUT(n1565) );
  INVX4 U736 ( .IN(C1_DATA7_2), .OUT(n987) );
  INVX4 U737 ( .IN(n879), .OUT(n692) );
  NANDX2 U738 ( .IN1(n429), .IN2(n903), .OUT(n879) );
  INVX4 U739 ( .IN(n651), .OUT(n865) );
  NANDX2 U740 ( .IN1(n650), .IN2(n649), .OUT(n651) );
  NANDX2 U741 ( .IN1(n1519), .IN2(n866), .OUT(n658) );
  NANDX2 U742 ( .IN1(n534), .IN2(n533), .OUT(n644) );
  INVX4 U743 ( .IN(n528), .OUT(n646) );
  NANDX2 U744 ( .IN1(n549), .IN2(n1298), .OUT(n890) );
  INVX4 U745 ( .IN(n582), .OUT(n615) );
  INVX4 U746 ( .IN(n558), .OUT(n559) );
  INVX4 U747 ( .IN(n536), .OUT(n537) );
  INVX4 U748 ( .IN(n548), .OUT(n908) );
  NANDX2 U749 ( .IN1(n504), .IN2(n505), .OUT(n641) );
  INVX4 U750 ( .IN(n499), .OUT(n670) );
  NANDX2 U751 ( .IN1(n639), .IN2(n868), .OUT(n905) );
  INVX4 U752 ( .IN(n556), .OUT(n673) );
  NANDX2 U753 ( .IN1(n485), .IN2(n868), .OUT(n486) );
  INVX4 U754 ( .IN(n484), .OUT(n868) );
  INVX4 U755 ( .IN(n639), .OUT(n485) );
  NANDX2 U756 ( .IN1(n469), .IN2(n1232), .OUT(n639) );
  INVX4 U757 ( .IN(n880), .OUT(n680) );
  NANDX2 U758 ( .IN1(n1484), .IN2(n503), .OUT(n880) );
  INVX4 U759 ( .IN(n501), .OUT(n667) );
  INVX4 U760 ( .IN(n502), .OUT(n1484) );
  NANDX2 U761 ( .IN1(n502), .IN2(n503), .OUT(n556) );
  INVX4 U762 ( .IN(n1510), .OUT(n503) );
  NANDX2 U763 ( .IN1(n1232), .IN2(n498), .OUT(n1510) );
  NANDX2 U764 ( .IN1(n1232), .IN2(n494), .OUT(n502) );
  INVX4 U765 ( .IN(n1505), .OUT(n1228) );
  NANDX2 U766 ( .IN1(n855), .IN2(n886), .OUT(n858) );
  NANDX2 U767 ( .IN1(n564), .IN2(n563), .OUT(n886) );
  INVX4 U768 ( .IN(n532), .OUT(n884) );
  NANDX2 U769 ( .IN1(n531), .IN2(n530), .OUT(n532) );
  INVX4 U770 ( .IN(n648), .OUT(n610) );
  INVX4 U771 ( .IN(n1498), .OUT(n530) );
  INVX4 U772 ( .IN(n529), .OUT(n645) );
  INVX4 U773 ( .IN(n1482), .OUT(n531) );
  INVX4 U774 ( .IN(n689), .OUT(n855) );
  NANDX2 U775 ( .IN1(n866), .IN2(n525), .OUT(n689) );
  INVX4 U776 ( .IN(n621), .OUT(n866) );
  INVX4 U777 ( .IN(n539), .OUT(n889) );
  INVX4 U778 ( .IN(n1290), .OUT(n1568) );
  INVX4 U779 ( .IN(n909), .OUT(n1298) );
  NANDX2 U780 ( .IN1(n430), .IN2(n698), .OUT(n697) );
  INVX1 U781 ( .IN(Adder_ack), .OUT(n430) );
  INVX4 U782 ( .IN(n875), .OUT(n897) );
  NANDX2 U783 ( .IN1(n1308), .IN2(n911), .OUT(n876) );
  NAND2X1 U784 ( .IN1(StateMC[1]), .IN2(n313), .OUT(n1606) );
  NAND2X1 U785 ( .IN1(StateMC[2]), .IN2(n300), .OUT(n550) );
  INVX4 U786 ( .IN(DP_OP_983_177_8739_n29), .OUT(DP_OP_983_177_8739_n11) );
  NANDX2 U787 ( .IN1(n199), .IN2(DP_OP_983_177_8739_n15), .OUT(
        DP_OP_983_177_8739_n29) );
  NANDX2 U788 ( .IN1(n199), .IN2(DP_OP_988_182_8739_n15), .OUT(
        DP_OP_988_182_8739_n25) );
  INVX4 U789 ( .IN(DP_OP_988_182_8739_n26), .OUT(DP_OP_988_182_8739_n15) );
  NANDX2 U790 ( .IN1(n207), .IN2(DP_OP_988_182_8739_n19), .OUT(
        DP_OP_988_182_8739_n26) );
  NANDX2 U791 ( .IN1(n199), .IN2(DP_OP_987_181_8739_n15), .OUT(
        DP_OP_987_181_8739_n29) );
  INVX4 U792 ( .IN(DP_OP_987_181_8739_n30), .OUT(DP_OP_987_181_8739_n15) );
  NANDX2 U793 ( .IN1(n207), .IN2(DP_OP_987_181_8739_n19), .OUT(
        DP_OP_987_181_8739_n30) );
  NANDX2 U794 ( .IN1(n199), .IN2(DP_OP_981_175_8739_n15), .OUT(
        DP_OP_981_175_8739_n29) );
  INVX4 U795 ( .IN(DP_OP_981_175_8739_n30), .OUT(DP_OP_981_175_8739_n15) );
  NANDX2 U796 ( .IN1(n207), .IN2(n369), .OUT(DP_OP_981_175_8739_n30) );
  NANDX2 U797 ( .IN1(n207), .IN2(DP_OP_984_178_8739_n19), .OUT(
        DP_OP_984_178_8739_n26) );
  NANDX2 U798 ( .IN1(n207), .IN2(DP_OP_985_179_8739_n19), .OUT(
        DP_OP_985_179_8739_n30) );
  NAND2X1 U799 ( .IN1(Datain1[12]), .IN2(n197), .OUT(n1136) );
  INVX4 U800 ( .IN(C1_DATA7_1), .OUT(n1139) );
  NANDX2 U801 ( .IN1(n1041), .IN2(n1040), .OUT(n1042) );
  NANDX2 U802 ( .IN1(n1041), .IN2(n1038), .OUT(n1039) );
  INVX4 U803 ( .IN(n1037), .OUT(n1038) );
  NANDX2 U804 ( .IN1(n396), .IN2(N2921), .OUT(n395) );
  INVX4 U805 ( .IN(n398), .OUT(DP_OP_979_173_2805_n58) );
  NANDX2 U806 ( .IN1(n396), .IN2(N2923), .OUT(n398) );
  INVX4 U807 ( .IN(n921), .OUT(N2923) );
  INVX4 U808 ( .IN(n1032), .OUT(n1197) );
  INVX4 U809 ( .IN(n1018), .OUT(n1191) );
  NANDX2 U810 ( .IN1(n1012), .IN2(n1503), .OUT(n1026) );
  INVX4 U811 ( .IN(n1010), .OUT(n1192) );
  NANDX2 U812 ( .IN1(n524), .IN2(n935), .OUT(n1008) );
  NANDX2 U813 ( .IN1(n476), .IN2(n482), .OUT(n1226) );
  INVX4 U814 ( .IN(n1007), .OUT(n1189) );
  NANDX2 U815 ( .IN1(n1203), .IN2(n1006), .OUT(n1007) );
  NANDX2 U816 ( .IN1(n483), .IN2(n482), .OUT(n1505) );
  INVX4 U817 ( .IN(n366), .OUT(n482) );
  INVX4 U818 ( .IN(n959), .OUT(n557) );
  INVX4 U819 ( .IN(n1004), .OUT(n1190) );
  NANDX2 U820 ( .IN1(n996), .IN2(n351), .OUT(n1187) );
  NANDX2 U821 ( .IN1(n492), .IN2(n1243), .OUT(n1027) );
  INVX4 U822 ( .IN(DP_OP_981_175_8739_n31), .OUT(n369) );
  INVX4 U823 ( .IN(DP_OP_981_175_8739_n32), .OUT(DP_OP_981_175_8739_n23) );
  NANDX2 U824 ( .IN1(n293), .IN2(DP_OP_985_179_8739_n27), .OUT(
        DP_OP_981_175_8739_n32) );
  INVX4 U825 ( .IN(n993), .OUT(n1188) );
  INVX4 U826 ( .IN(n985), .OUT(n1181) );
  INVX4 U827 ( .IN(DP_OP_984_178_8739_n27), .OUT(DP_OP_984_178_8739_n19) );
  INVX4 U828 ( .IN(n978), .OUT(n1271) );
  INVX4 U829 ( .IN(DP_OP_985_179_8739_n31), .OUT(DP_OP_985_179_8739_n19) );
  NANDX2 U830 ( .IN1(n975), .IN2(n974), .OUT(n1184) );
  NANDX2 U831 ( .IN1(n979), .IN2(n1306), .OUT(n1499) );
  NANDX2 U832 ( .IN1(n468), .IN2(n467), .OUT(n1232) );
  INVX4 U833 ( .IN(n466), .OUT(n467) );
  NANDX2 U834 ( .IN1(n1011), .IN2(n1233), .OUT(n466) );
  NANDX2 U835 ( .IN1(n460), .IN2(n1523), .OUT(n1233) );
  NANDX2 U836 ( .IN1(n459), .IN2(n1523), .OUT(n1011) );
  INVX4 U837 ( .IN(n954), .OUT(n1523) );
  INVX4 U838 ( .IN(n455), .OUT(n669) );
  INVX4 U839 ( .IN(n414), .OUT(n1485) );
  NANDX2 U840 ( .IN1(n671), .IN2(n1501), .OUT(n1243) );
  INVX4 U841 ( .IN(n904), .OUT(n1501) );
  NANDX2 U842 ( .IN1(n224), .IN2(n490), .OUT(n904) );
  NANDX2 U843 ( .IN1(n481), .IN2(n520), .OUT(n959) );
  NANDX2 U844 ( .IN1(n480), .IN2(n479), .OUT(n958) );
  INVX4 U845 ( .IN(n475), .OUT(n965) );
  NANDX2 U846 ( .IN1(n379), .IN2(n474), .OUT(n475) );
  INVX4 U847 ( .IN(n950), .OUT(n623) );
  NANDX2 U848 ( .IN1(n454), .IN2(n458), .OUT(n1500) );
  NANDX2 U849 ( .IN1(n490), .IN2(n458), .OUT(n954) );
  INVX4 U850 ( .IN(n472), .OUT(n458) );
  NANDX2 U851 ( .IN1(n453), .IN2(n600), .OUT(n472) );
  NANDX2 U852 ( .IN1(n373), .IN2(n372), .OUT(n600) );
  INVX4 U853 ( .IN(n896), .OUT(n490) );
  NANDX2 U854 ( .IN1(n336), .IN2(n489), .OUT(n896) );
  NANDX2 U855 ( .IN1(n450), .IN2(n487), .OUT(n451) );
  INVX4 U856 ( .IN(n491), .OUT(n487) );
  NANDX2 U857 ( .IN1(n358), .IN2(n449), .OUT(n491) );
  INVX4 U858 ( .IN(n359), .OUT(n358) );
  NANDX2 U859 ( .IN1(n445), .IN2(n446), .OUT(n359) );
  NANDX2 U860 ( .IN1(n1211), .IN2(n953), .OUT(n955) );
  INVX4 U861 ( .IN(n471), .OUT(n686) );
  NANDX2 U862 ( .IN1(n331), .IN2(n330), .OUT(n471) );
  INVX4 U863 ( .IN(n360), .OUT(n445) );
  NANDX2 U864 ( .IN1(n463), .IN2(n462), .OUT(n500) );
  NANDX2 U865 ( .IN1(n329), .IN2(n477), .OUT(n462) );
  INVX4 U866 ( .IN(n478), .OUT(n477) );
  NANDX2 U867 ( .IN1(n297), .IN2(n299), .OUT(n478) );
  NANDX2 U868 ( .IN1(n949), .IN2(n948), .OUT(n998) );
  INVX4 U869 ( .IN(n947), .OUT(n949) );
  NANDX2 U870 ( .IN1(n1518), .IN2(n946), .OUT(n947) );
  INVX4 U871 ( .IN(n979), .OUT(n1518) );
  NANDX2 U872 ( .IN1(n538), .IN2(n507), .OUT(n979) );
  NANDX2 U873 ( .IN1(n997), .IN2(n943), .OUT(n1037) );
  NANDX2 U874 ( .IN1(n941), .IN2(n1211), .OUT(n946) );
  INVX4 U875 ( .IN(n1235), .OUT(n1211) );
  NANDX2 U876 ( .IN1(n516), .IN2(n1520), .OUT(n1212) );
  NANDX2 U877 ( .IN1(n514), .IN2(n1520), .OUT(n1487) );
  NANDX2 U878 ( .IN1(n1000), .IN2(n1239), .OUT(n1210) );
  INVX4 U879 ( .IN(n1492), .OUT(n1000) );
  INVX4 U880 ( .IN(n940), .OUT(n948) );
  INVX4 U881 ( .IN(n1251), .OUT(n975) );
  NANDX2 U882 ( .IN1(n419), .IN2(n521), .OUT(n936) );
  NANDX2 U883 ( .IN1(n932), .IN2(n1279), .OUT(n1203) );
  INVX4 U884 ( .IN(n1227), .OUT(n1279) );
  NANDX2 U885 ( .IN1(n931), .IN2(n930), .OUT(n1227) );
  INVX4 U886 ( .IN(n523), .OUT(n935) );
  NANDX2 U887 ( .IN1(n522), .IN2(n521), .OUT(n523) );
  INVX4 U888 ( .IN(n1491), .OUT(n1205) );
  NANDX2 U889 ( .IN1(n519), .IN2(n521), .OUT(n1491) );
  INVX4 U890 ( .IN(n513), .OUT(n521) );
  NANDX2 U891 ( .IN1(n512), .IN2(n1520), .OUT(n513) );
  INVX4 U892 ( .IN(n511), .OUT(n1520) );
  NANDX2 U893 ( .IN1(n510), .IN2(n1488), .OUT(n511) );
  NANDX2 U894 ( .IN1(n1214), .IN2(n995), .OUT(n997) );
  INVX4 U895 ( .IN(n1246), .OUT(n995) );
  NANDX2 U896 ( .IN1(n929), .IN2(n1244), .OUT(n1246) );
  INVX4 U897 ( .IN(n928), .OUT(n1214) );
  NANDX2 U898 ( .IN1(n1216), .IN2(n1244), .OUT(n1041) );
  INVX4 U899 ( .IN(n927), .OUT(n1216) );
  INVX4 U900 ( .IN(n509), .OUT(n1488) );
  NANDX2 U901 ( .IN1(n409), .IN2(n210), .OUT(n397) );
  NANDX2 U902 ( .IN1(DP_OP_979_173_2805_n52), .IN2(DP_OP_990_184_2805_n58), 
        .OUT(DP_OP_990_184_2805_n51) );
  NANDX2 U903 ( .IN1(n918), .IN2(n1237), .OUT(n919) );
  NANDX2 U904 ( .IN1(n210), .IN2(n1230), .OUT(n1244) );
  INVX4 U905 ( .IN(n992), .OUT(n1230) );
  INVX4 U906 ( .IN(n917), .OUT(n930) );
  INVX4 U907 ( .IN(n1219), .OUT(n918) );
  NANDX2 U908 ( .IN1(Final_Mantissa_reg[10]), .IN2(n538), .OUT(n506) );
  NANDX2 U909 ( .IN1(n923), .IN2(n976), .OUT(n1257) );
  INVX4 U910 ( .IN(n1494), .OUT(n976) );
  NANDX2 U911 ( .IN1(n1548), .IN2(n1502), .OUT(n1494) );
  INVX4 U912 ( .IN(n977), .OUT(n923) );
  INVX4 U913 ( .IN(DP_OP_979_173_2805_n76), .OUT(n409) );
  NANDX2 U914 ( .IN1(n1387), .IN2(n197), .OUT(n1462) );
  INVX4 U915 ( .IN(n1421), .OUT(n1351) );
  NANDX2 U916 ( .IN1(n418), .IN2(n1427), .OUT(n1348) );
  INVX4 U917 ( .IN(n1467), .OUT(n1456) );
  NANDX2 U918 ( .IN1(n376), .IN2(n378), .OUT(n1467) );
  INVX4 U919 ( .IN(n377), .OUT(n376) );
  NANDX2 U920 ( .IN1(n1411), .IN2(n1406), .OUT(n377) );
  INVX4 U921 ( .IN(n1426), .OUT(n1451) );
  NANDX2 U922 ( .IN1(n1345), .IN2(n1384), .OUT(n1426) );
  INVX4 U923 ( .IN(n1323), .OUT(n1427) );
  NANDX2 U924 ( .IN1(n1357), .IN2(n1443), .OUT(n1421) );
  INVX4 U925 ( .IN(n748), .OUT(n1357) );
  INVX4 U926 ( .IN(N147), .OUT(n769) );
  NANDX2 U927 ( .IN1(n1406), .IN2(n378), .OUT(n375) );
  INVX4 U928 ( .IN(n1425), .OUT(n1409) );
  NANDX2 U929 ( .IN1(n382), .IN2(n378), .OUT(n1425) );
  NANDX2 U930 ( .IN1(n1345), .IN2(n1405), .OUT(n794) );
  INVX4 U931 ( .IN(n1398), .OUT(n1402) );
  NANDX2 U932 ( .IN1(n1397), .IN2(n1443), .OUT(n1453) );
  NANDX2 U933 ( .IN1(n1332), .IN2(n1620), .OUT(n1387) );
  INVX4 U934 ( .IN(n1408), .OUT(n1386) );
  INVX4 U935 ( .IN(n1320), .OUT(n1384) );
  NANDX2 U936 ( .IN1(n400), .IN2(n722), .OUT(n399) );
  INVX4 U937 ( .IN(n401), .OUT(n400) );
  INVX4 U938 ( .IN(n388), .OUT(n345) );
  INVX4 U939 ( .IN(n1383), .OUT(n1385) );
  NANDX2 U940 ( .IN1(n1382), .IN2(n1381), .OUT(n1383) );
  NANDX2 U941 ( .IN1(n198), .IN2(n1345), .OUT(n1369) );
  BUF4X U942 ( .IN(Datain1[6]), .OUT(n418) );
  BUF4X U943 ( .IN(Datain1[5]), .OUT(n417) );
  BUF4X U944 ( .IN(Datain1[4]), .OUT(n416) );
  NANDX2 U945 ( .IN1(n198), .IN2(N419), .OUT(n1350) );
  INVX4 U946 ( .IN(n1627), .OUT(n1534) );
  NANDX2 U947 ( .IN1(n753), .IN2(n1401), .OUT(n772) );
  INVX4 U948 ( .IN(n752), .OUT(n1401) );
  NANDX2 U949 ( .IN1(n390), .IN2(n389), .OUT(n385) );
  NANDX2 U950 ( .IN1(n1603), .IN2(n1602), .OUT(n389) );
  BUF4X U951 ( .IN(Datain2[12]), .OUT(DP_OP_982J1_125_6202_n180) );
  NAND2X1 U952 ( .IN1(Datain1[13]), .IN2(n1604), .OUT(n392) );
  BUF4X U953 ( .IN(Datain2[13]), .OUT(DP_OP_982J1_125_6202_n181) );
  BUF4X U954 ( .IN(Datain2[7]), .OUT(DP_OP_982J1_125_6202_n175) );
  NANDX2 U955 ( .IN1(n1591), .IN2(Data_valid), .OUT(n1605) );
  NAND2X1 U956 ( .IN1(n300), .IN2(n313), .OUT(n1580) );
  NAND2X1 U957 ( .IN1(Adder_ack), .IN2(n698), .OUT(n1290) );
  NAND2X1 U958 ( .IN1(n225), .IN2(n197), .OUT(n1119) );
  INVX4 U959 ( .IN(n294), .OUT(DP_OP_979_173_2805_n76) );
  NAND2X1 U960 ( .IN1(n1556), .IN2(n1551), .OUT(n1480) );
  NAND2X1 U961 ( .IN1(n1556), .IN2(n1561), .OUT(n1543) );
  INVX1 U962 ( .IN(n1625), .OUT(n1557) );
  NAND2X1 U963 ( .IN1(n429), .IN2(n307), .OUT(n1310) );
  NAND2X1 U964 ( .IN1(n1556), .IN2(n1306), .OUT(n1307) );
  NAND2X1 U965 ( .IN1(n429), .IN2(n909), .OUT(n910) );
  NAND2X1 U966 ( .IN1(add_x_35_A_4_), .IN2(add_x_35_A_5_), .OUT(n1540) );
  INVX1 U967 ( .IN(n1536), .OUT(n112) );
  INVX1 U968 ( .IN(n1528), .OUT(n111) );
  NAND2X1 U969 ( .IN1(n1523), .IN2(n1522), .OUT(n1524) );
  INVX1 U970 ( .IN(n1515), .OUT(n110) );
  NAND2X1 U971 ( .IN1(n1521), .IN2(n1493), .OUT(n1495) );
  INVX1 U972 ( .IN(Exc_Ack), .OUT(n1259) );
  NAND2X1 U973 ( .IN1(Final_Mantissa_reg[10]), .IN2(n890), .OUT(n899) );
  INVX1 U974 ( .IN(n1519), .OUT(n885) );
  INVX1 U975 ( .IN(n793), .OUT(n796) );
  NAND2X1 U976 ( .IN1(N160), .IN2(N161), .OUT(n777) );
  INVX1 U977 ( .IN(N160), .OUT(n773) );
  INVX1 U978 ( .IN(N149), .OUT(n763) );
  NAND2X1 U979 ( .IN1(N148), .IN2(N149), .OUT(n765) );
  NAND2X1 U980 ( .IN1(Exc_Ack), .IN2(n415), .OUT(n1577) );
  INVX1 U981 ( .IN(n1225), .OUT(n1256) );
  NAND2X1 U982 ( .IN1(n1494), .IN2(n1274), .OUT(n1483) );
  INVX1 U983 ( .IN(n1237), .OUT(n1240) );
  INVX1 U984 ( .IN(n1233), .OUT(n1236) );
  INVX1 U985 ( .IN(n1232), .OUT(n1252) );
  INVX1 U986 ( .IN(n1506), .OUT(n1231) );
  INVX1 U987 ( .IN(n1487), .OUT(n1217) );
  INVX1 U988 ( .IN(C1_DATA7_7), .OUT(n1183) );
  NAND2X1 U989 ( .IN1(Datain1[0]), .IN2(n1456), .OUT(n1340) );
  INVX1 U990 ( .IN(n1462), .OUT(n1396) );
  NAND2X1 U991 ( .IN1(n202), .IN2(n1358), .OUT(n1326) );
  INVX1 U992 ( .IN(n1175), .OUT(n1176) );
  NAND2X1 U993 ( .IN1(n341), .IN2(DP_OP_990_184_2805_n13), .OUT(n340) );
  NAND2X1 U994 ( .IN1(DP_OP_979_173_2805_n77), .IN2(DP_OP_990_184_2805_n14), 
        .OUT(n341) );
  NAND2X1 U995 ( .IN1(N144), .IN2(N145), .OUT(n829) );
  INVX1 U996 ( .IN(N145), .OUT(n826) );
  INVX1 U997 ( .IN(n825), .OUT(n849) );
  INVX1 U998 ( .IN(n821), .OUT(n822) );
  NAND2X1 U999 ( .IN1(N156), .IN2(N157), .OUT(n805) );
  INVX1 U1000 ( .IN(N157), .OUT(n803) );
  NAND2X1 U1001 ( .IN1(n423), .IN2(n615), .OUT(n614) );
  INVX1 U1002 ( .IN(n747), .OUT(n755) );
  INVX1 U1003 ( .IN(Datain2[2]), .OUT(n830) );
  NAND2X1 U1004 ( .IN1(N152), .IN2(N153), .OUT(n731) );
  INVX1 U1005 ( .IN(N153), .OUT(n729) );
  INVX1 U1006 ( .IN(Datain2[3]), .OUT(n827) );
  INVX1 U1007 ( .IN(N152), .OUT(n727) );
  INVX1 U1008 ( .IN(n721), .OUT(n724) );
  INVX1 U1009 ( .IN(Datain1[2]), .OUT(n1312) );
  NAND2X1 U1010 ( .IN1(N164), .IN2(N165), .OUT(n705) );
  INVX1 U1011 ( .IN(N165), .OUT(n703) );
  NAND2X1 U1012 ( .IN1(n1260), .IN2(n702), .OUT(n802) );
  INVX1 U1013 ( .IN(n698), .OUT(n700) );
  NAND2X1 U1014 ( .IN1(StateMC[1]), .IN2(n1566), .OUT(n1297) );
  BUF4X U1015 ( .IN(n1567), .OUT(n415) );
  NAND2X1 U1016 ( .IN1(n1197), .IN2(C1_DATA1_2), .OUT(n1033) );
  INVX1 U1017 ( .IN(n600), .OUT(n668) );
  NAND2X1 U1018 ( .IN1(n897), .IN2(n221), .OUT(n653) );
  NAND2X1 U1019 ( .IN1(n308), .IN2(n477), .OUT(n535) );
  NAND2X1 U1020 ( .IN1(n502), .IN2(n1510), .OUT(n499) );
  NAND2X1 U1021 ( .IN1(n856), .IN2(n903), .OUT(n857) );
  NAND2X1 U1022 ( .IN1(n426), .IN2(n645), .OUT(n564) );
  INVX1 U1023 ( .IN(n1606), .OUT(n551) );
  INVX1 U1024 ( .IN(n1134), .OUT(n1135) );
  NAND2X1 U1025 ( .IN1(n1197), .IN2(C1_DATA1_5), .OUT(n1128) );
  INVX1 U1026 ( .IN(n1151), .OUT(n1152) );
  INVX1 U1027 ( .IN(n1117), .OUT(n1118) );
  INVX1 U1028 ( .IN(n1234), .OUT(n1012) );
  NAND2X1 U1029 ( .IN1(n1499), .IN2(n1201), .OUT(n1009) );
  NAND2X1 U1030 ( .IN1(n1499), .IN2(n1204), .OUT(n1005) );
  INVX1 U1031 ( .IN(DP_OP_982_176_8739_n23), .OUT(DP_OP_982_176_8739_n19) );
  NAND2X1 U1032 ( .IN1(n409), .IN2(n293), .OUT(DP_OP_982_176_8739_n23) );
  NAND2X1 U1033 ( .IN1(n998), .IN2(n994), .OUT(n352) );
  INVX1 U1034 ( .IN(n1027), .OUT(n1247) );
  NAND2X1 U1035 ( .IN1(n992), .IN2(n990), .OUT(n993) );
  NAND2X1 U1036 ( .IN1(n1205), .IN2(n1499), .OUT(n989) );
  INVX1 U1037 ( .IN(n958), .OUT(n365) );
  NAND2X1 U1038 ( .IN1(n1202), .IN2(n1499), .OUT(n973) );
  INVX1 U1039 ( .IN(n1521), .OUT(n1306) );
  INVX1 U1040 ( .IN(n1023), .OUT(n967) );
  NAND2X1 U1041 ( .IN1(n1244), .IN2(n966), .OUT(n1023) );
  INVX1 U1042 ( .IN(n1243), .OUT(n966) );
  NAND2X1 U1043 ( .IN1(n959), .IN2(n1203), .OUT(n960) );
  NAND2X1 U1044 ( .IN1(n427), .IN2(n297), .OUT(n481) );
  NAND2X1 U1045 ( .IN1(n312), .IN2(n478), .OUT(n479) );
  INVX1 U1046 ( .IN(n1014), .OUT(n957) );
  NAND2X1 U1047 ( .IN1(n309), .IN2(n186), .OUT(n374) );
  INVX1 U1048 ( .IN(n952), .OUT(n953) );
  NAND2X1 U1049 ( .IN1(n1492), .IN2(n394), .OUT(n945) );
  NAND2X1 U1050 ( .IN1(n1492), .IN2(n1521), .OUT(n393) );
  NAND2X1 U1051 ( .IN1(n292), .IN2(n1230), .OUT(n937) );
  NAND2X1 U1052 ( .IN1(n292), .IN2(n1239), .OUT(n929) );
  INVX1 U1053 ( .IN(n397), .OUT(DP_OP_980_174_8739_n19) );
  BUF4X U1054 ( .IN(Final_Exponent_reg[1]), .OUT(n407) );
  INVX1 U1055 ( .IN(n538), .OUT(n1502) );
  INVX4 U1056 ( .IN(n408), .OUT(DP_OP_979_173_2805_n77) );
  INVX4 U1057 ( .IN(n304), .OUT(DP_OP_979_173_2805_n78) );
  INVX4 U1058 ( .IN(n295), .OUT(DP_OP_979_173_2805_n79) );
  INVX1 U1059 ( .IN(Datain1[3]), .OUT(n1321) );
  INVX1 U1060 ( .IN(Datain1[1]), .OUT(n1322) );
  INVX1 U1061 ( .IN(n1353), .OUT(n1354) );
  NAND2X1 U1062 ( .IN1(Datain2[5]), .IN2(n1397), .OUT(n1353) );
  NAND2X1 U1063 ( .IN1(n1395), .IN2(n1351), .OUT(n1365) );
  INVX1 U1064 ( .IN(n1370), .OUT(n1347) );
  INVX1 U1065 ( .IN(Datain2[4]), .OUT(n1330) );
  NAND2X1 U1066 ( .IN1(N362), .IN2(n1424), .OUT(n1414) );
  NAND2X1 U1067 ( .IN1(N364), .IN2(n1397), .OUT(n357) );
  NAND2X1 U1068 ( .IN1(Datain2[3]), .IN2(n197), .OUT(n1404) );
  NAND2X1 U1069 ( .IN1(N364), .IN2(n1401), .OUT(n1361) );
  INVX1 U1070 ( .IN(Datain2[6]), .OUT(n1352) );
  INVX1 U1071 ( .IN(n1417), .OUT(n1375) );
  INVX1 U1072 ( .IN(N364), .OUT(n753) );
  INVX1 U1073 ( .IN(n434), .OUT(n387) );
  INVX4 U1074 ( .IN(n293), .OUT(n411) );
  BUF4X U1075 ( .IN(Final_Mantissa_reg[4]), .OUT(n420) );
  BUF4X U1076 ( .IN(Final_Mantissa_reg[3]), .OUT(n419) );
  BUF4X U1077 ( .IN(Final_Mantissa_reg[9]), .OUT(n424) );
  INVX1 U1078 ( .IN(DP_OP_983_177_8739_n15), .OUT(DP_OP_983_177_8739_n30) );
  INVX1 U1079 ( .IN(n946), .OUT(n984) );
  NAND2X1 U1080 ( .IN1(n386), .IN2(n385), .OUT(n384) );
  BUF4X U1081 ( .IN(Final_Mantissa_reg[8]), .OUT(n425) );
  MUX2X1 U1082 ( .IN1(n327), .IN2(n326), .S(n325), .OUT(n404) );
  OAI21 U1083 ( .IN1(n333), .IN2(n478), .IN3(n420), .OUT(n330) );
  NOR2X1 U1084 ( .IN1(n420), .IN2(n333), .OUT(n332) );
  NOR2X1 U1085 ( .IN1(n455), .IN2(n896), .OUT(n454) );
  AOI21 U1086 ( .IN1(n342), .IN2(n339), .IN3(n1627), .OUT(n1175) );
  NOR2X1 U1087 ( .IN1(n1172), .IN2(n343), .OUT(n342) );
  AOI21 U1088 ( .IN1(n1186), .IN2(C1_DATA2_4), .IN3(n1168), .OUT(n344) );
  INVX4 U1089 ( .IN(n399), .OUT(n1405) );
  NANDX2 U1090 ( .IN1(n438), .IN2(n345), .OUT(n1318) );
  OAI21 U1091 ( .IN1(n349), .IN2(n348), .IN3(n1534), .OUT(n347) );
  NAND3X1 U1092 ( .IN1(n364), .IN2(n1500), .IN3(n965), .OUT(n363) );
  NAND3X1 U1093 ( .IN1(n958), .IN2(n965), .IN3(n1500), .OUT(n1506) );
  NOR2X1 U1094 ( .IN1(n365), .IN2(n1485), .OUT(n364) );
  AOI22 U1095 ( .IN1(n680), .IN2(n959), .IN3(n426), .IN4(n673), .OUT(n638) );
  OAI21 U1096 ( .IN1(n368), .IN2(n794), .IN3(n1564), .OUT(n723) );
  NOR2X1 U1097 ( .IN1(n198), .IN2(n1411), .OUT(n368) );
  OAI21 U1098 ( .IN1(n374), .IN2(n457), .IN3(n371), .OUT(n370) );
  INVX4 U1099 ( .IN(n794), .OUT(n378) );
  INVX4 U1100 ( .IN(n375), .OUT(n1446) );
  NOR2X1 U1101 ( .IN1(DP_OP_979_173_2805_n77), .IN2(DP_OP_982_176_8739_n23), 
        .OUT(DP_OP_982_176_8739_n15) );
  MUX2X1 U1102 ( .IN1(n1340), .IN2(n1371), .S(n202), .OUT(n1341) );
  NANDX2 U1103 ( .IN1(n434), .IN2(n385), .OUT(n1388) );
  NOR2X1 U1104 ( .IN1(n387), .IN2(N362), .OUT(n386) );
  INVX1 U1105 ( .IN(n1017), .OUT(n394) );
  OAI21 U1106 ( .IN1(n404), .IN2(n825), .IN3(n402), .OUT(n1070) );
  INVX4 U1107 ( .IN(n405), .OUT(DP_OP_979_173_2805_n80) );
  TIEHI U1108 ( .OUT(n73) );
  INVX1 U1109 ( .IN(DP_OP_981_175_8739_n7), .OUT(DP_OP_981_175_8739_n28) );
  INVX1 U1110 ( .IN(DP_OP_983_177_8739_n19), .OUT(DP_OP_983_177_8739_n31) );
  NOR2X1 U1111 ( .IN1(n384), .IN2(n772), .OUT(n412) );
  INVX1 U1112 ( .IN(N161), .OUT(n775) );
  NAND2X1 U1113 ( .IN1(Datain1[9]), .IN2(n197), .OUT(n1046) );
  NAND2X1 U1114 ( .IN1(Datain1[8]), .IN2(n197), .OUT(n1153) );
  NOR2X1 U1115 ( .IN1(StateMC[0]), .IN2(n313), .OUT(n1566) );
  INVX4 U1116 ( .IN(n1581), .OUT(n901) );
  NANDX2 U1117 ( .IN1(n429), .IN2(n901), .OUT(n1627) );
  NOR2X1 U1118 ( .IN1(n301), .IN2(n1606), .OUT(n698) );
  NOR2X1 U1119 ( .IN1(RSTn_BAR), .IN2(n1290), .OUT(n913) );
  NOR2X1 U1120 ( .IN1(StateMC[0]), .IN2(n1606), .OUT(n1626) );
  AOI21 U1121 ( .IN1(n1298), .IN2(n551), .IN3(n1310), .OUT(n432) );
  AOI21 U1122 ( .IN1(Adder_dataout[8]), .IN2(n913), .IN3(n432), .OUT(n433) );
  NOR2X1 U1123 ( .IN1(RSTn_BAR), .IN2(n1605), .OUT(n434) );
  NOR2X1 U1124 ( .IN1(StateMC[1]), .IN2(StateMC[0]), .OUT(n435) );
  AOI21 U1125 ( .IN1(n1592), .IN2(n435), .IN3(RSTn_BAR), .OUT(n924) );
  NOR2X1 U1126 ( .IN1(n1534), .IN2(n924), .OUT(n1622) );
  INVX4 U1127 ( .IN(n413), .OUT(n1465) );
  NOR2X1 U1128 ( .IN1(n437), .IN2(n1605), .OUT(n438) );
  AOI22 U1129 ( .IN1(Op2_Sign_reg), .IN2(n1465), .IN3(Datain1[15]), .IN4(n1564), .OUT(n439) );
  OAI21 U1130 ( .IN1(n1388), .IN2(n440), .IN3(n439), .OUT(n1090) );
  AOI22 U1131 ( .IN1(Op1_Sign_reg), .IN2(n1465), .IN3(Datain2[15]), .IN4(n1564), .OUT(n441) );
  OAI21 U1132 ( .IN1(n1388), .IN2(n442), .IN3(n441), .OUT(n1081) );
  NOR2X1 U1133 ( .IN1(n426), .IN2(n421), .OUT(n444) );
  NAND3X1 U1134 ( .IN1(n444), .IN2(n445), .IN3(n443), .OUT(n457) );
  MUX2X1 U1135 ( .IN1(n186), .IN2(n422), .S(n457), .OUT(n455) );
  NOR2X1 U1136 ( .IN1(n425), .IN2(n424), .OUT(n450) );
  NOR2X1 U1137 ( .IN1(n423), .IN2(n421), .OUT(n446) );
  NOR2X1 U1138 ( .IN1(n448), .IN2(n447), .OUT(n449) );
  NAND3X1 U1139 ( .IN1(n425), .IN2(n424), .IN3(n491), .OUT(n452) );
  OAI21 U1140 ( .IN1(n420), .IN2(n462), .IN3(n421), .OUT(n456) );
  NOR2X1 U1141 ( .IN1(n669), .IN2(n950), .OUT(n459) );
  NOR2X1 U1142 ( .IN1(n669), .IN2(n952), .OUT(n460) );
  NAND3X1 U1143 ( .IN1(n1500), .IN2(n1011), .IN3(n1233), .OUT(n461) );
  OAI21 U1144 ( .IN1(n428), .IN2(n478), .IN3(n419), .OUT(n463) );
  NOR2X1 U1145 ( .IN1(n500), .IN2(n954), .OUT(n464) );
  NOR2X1 U1146 ( .IN1(carry_reg), .IN2(n508), .OUT(n1509) );
  NAND3X1 U1147 ( .IN1(n426), .IN2(n427), .IN3(n428), .OUT(n470) );
  NOR2X1 U1148 ( .IN1(n623), .IN2(n896), .OUT(n474) );
  NOR2X1 U1149 ( .IN1(n557), .IN2(n958), .OUT(n483) );
  NAND3X1 U1150 ( .IN1(n1226), .IN2(n1506), .IN3(n1505), .OUT(n577) );
  NOR2X1 U1151 ( .IN1(n1485), .IN2(n577), .OUT(n1522) );
  INVX4 U1152 ( .IN(n486), .OUT(n903) );
  NOR2X1 U1153 ( .IN1(n600), .IN2(n904), .OUT(n492) );
  MUX2X1 U1154 ( .IN1(n425), .IN2(n314), .S(n192), .OUT(n671) );
  NAND3X1 U1155 ( .IN1(n920), .IN2(n1027), .IN3(n1011), .OUT(n493) );
  NOR2X1 U1156 ( .IN1(n493), .IN2(n1228), .OUT(n494) );
  NAND3X1 U1157 ( .IN1(n1243), .IN2(n1027), .IN3(n1233), .OUT(n495) );
  AOI22 U1158 ( .IN1(n670), .IN2(n958), .IN3(n951), .IN4(n667), .OUT(n505) );
  AOI22 U1159 ( .IN1(n673), .IN2(n686), .IN3(n623), .IN4(n680), .OUT(n504) );
  INVX4 U1160 ( .IN(n1223), .OUT(n1272) );
  NOR2X1 U1161 ( .IN1(Final_Mantissa_reg[10]), .IN2(n1556), .OUT(n507) );
  NOR2X1 U1162 ( .IN1(n303), .IN2(n508), .OUT(n1521) );
  OAI21 U1163 ( .IN1(n1272), .IN2(n1499), .IN3(n901), .OUT(n621) );
  NOR2X1 U1164 ( .IN1(n420), .IN2(n515), .OUT(n512) );
  NOR2X1 U1165 ( .IN1(n425), .IN2(n423), .OUT(n510) );
  NOR2X1 U1166 ( .IN1(n422), .IN2(n311), .OUT(n514) );
  NOR2X1 U1167 ( .IN1(n298), .IN2(n515), .OUT(n516) );
  NAND3X1 U1168 ( .IN1(n1492), .IN2(n1487), .IN3(n1212), .OUT(n517) );
  NOR2X1 U1169 ( .IN1(n419), .IN2(n312), .OUT(n519) );
  NOR2X1 U1170 ( .IN1(n428), .IN2(n419), .OUT(n522) );
  NAND3X1 U1171 ( .IN1(n1491), .IN2(n1008), .IN3(n1493), .OUT(n864) );
  NOR2X1 U1172 ( .IN1(n1519), .IN2(n864), .OUT(n525) );
  AOI22 U1173 ( .IN1(n428), .IN2(n646), .IN3(n420), .IN4(n610), .OUT(n534) );
  AOI22 U1174 ( .IN1(n645), .IN2(n419), .IN3(n421), .IN4(n884), .OUT(n533) );
  AOI22 U1175 ( .IN1(n610), .IN2(n426), .IN3(n427), .IN4(n884), .OUT(n544) );
  NOR2X1 U1176 ( .IN1(n301), .IN2(n550), .OUT(n1563) );
  OAI21 U1177 ( .IN1(n421), .IN2(n537), .IN3(n558), .OUT(n541) );
  AOI22 U1178 ( .IN1(n1568), .IN2(Adder_dataout[2]), .IN3(n422), .IN4(n889), 
        .OUT(n540) );
  OAI21 U1179 ( .IN1(n893), .IN2(n541), .IN3(n540), .OUT(n542) );
  AOI21 U1180 ( .IN1(n623), .IN2(n897), .IN3(n542), .OUT(n543) );
  OAI21 U1181 ( .IN1(n658), .IN2(n544), .IN3(n543), .OUT(n545) );
  AOI21 U1182 ( .IN1(n855), .IN2(n644), .IN3(n545), .OUT(n546) );
  OAI21 U1183 ( .IN1(n905), .IN2(n638), .IN3(n546), .OUT(n547) );
  AOI21 U1184 ( .IN1(n903), .IN2(n641), .IN3(n547), .OUT(n554) );
  NOR2X1 U1185 ( .IN1(n551), .IN2(n1309), .OUT(n906) );
  OAI21 U1186 ( .IN1(RSTn_BAR), .IN2(n552), .IN3(n911), .OUT(n694) );
  OAI21 U1187 ( .IN1(RSTn_BAR), .IN2(n554), .IN3(n553), .OUT(n1067) );
  AOI22 U1188 ( .IN1(n667), .IN2(n426), .IN3(n680), .IN4(n958), .OUT(n555) );
  OAI21 U1189 ( .IN1(n557), .IN2(n556), .IN3(n555), .OUT(n856) );
  OAI21 U1190 ( .IN1(n422), .IN2(n559), .IN3(n582), .OUT(n561) );
  AOI22 U1191 ( .IN1(n1568), .IN2(Adder_dataout[3]), .IN3(n423), .IN4(n889), 
        .OUT(n560) );
  OAI21 U1192 ( .IN1(n893), .IN2(n561), .IN3(n560), .OUT(n562) );
  AOI21 U1193 ( .IN1(n897), .IN2(n669), .IN3(n562), .OUT(n570) );
  AOI22 U1194 ( .IN1(n610), .IN2(n427), .IN3(n428), .IN4(n884), .OUT(n563) );
  AOI22 U1195 ( .IN1(n645), .IN2(n420), .IN3(n422), .IN4(n884), .OUT(n566) );
  AOI22 U1196 ( .IN1(n419), .IN2(n646), .IN3(n421), .IN4(n610), .OUT(n565) );
  AOI21 U1197 ( .IN1(n566), .IN2(n565), .IN3(n689), .OUT(n567) );
  NAND3X1 U1198 ( .IN1(n570), .IN2(n569), .IN3(n568), .OUT(n571) );
  AOI21 U1199 ( .IN1(n679), .IN2(n856), .IN3(n571), .OUT(n576) );
  AOI22 U1200 ( .IN1(n951), .IN2(n670), .IN3(n686), .IN4(n667), .OUT(n573) );
  AOI22 U1201 ( .IN1(n673), .IN2(n623), .IN3(n680), .IN4(n669), .OUT(n572) );
  AOI22 U1202 ( .IN1(n422), .IN2(n694), .IN3(n574), .IN4(n692), .OUT(n575) );
  OAI21 U1203 ( .IN1(RSTn_BAR), .IN2(n576), .IN3(n575), .OUT(n1066) );
  NAND3X1 U1204 ( .IN1(n866), .IN2(n864), .IN3(n884), .OUT(n579) );
  OAI21 U1205 ( .IN1(n880), .IN2(n640), .IN3(n579), .OUT(n599) );
  AOI22 U1206 ( .IN1(n670), .IN2(n959), .IN3(n958), .IN4(n667), .OUT(n581) );
  AOI22 U1207 ( .IN1(n673), .IN2(n951), .IN3(n680), .IN4(n686), .OUT(n580) );
  AOI22 U1208 ( .IN1(n427), .IN2(n646), .IN3(n419), .IN4(n610), .OUT(n585) );
  AOI22 U1209 ( .IN1(n645), .IN2(n428), .IN3(n420), .IN4(n884), .OUT(n584) );
  AOI22 U1210 ( .IN1(n646), .IN2(n421), .IN3(n422), .IN4(n645), .OUT(n587) );
  OAI21 U1211 ( .IN1(n309), .IN2(n648), .IN3(n587), .OUT(n593) );
  AOI22 U1212 ( .IN1(n1568), .IN2(Adder_dataout[5]), .IN3(n424), .IN4(n889), 
        .OUT(n588) );
  AOI21 U1213 ( .IN1(n897), .IN2(n671), .IN3(n589), .OUT(n590) );
  OAI21 U1214 ( .IN1(n591), .IN2(n614), .IN3(n590), .OUT(n592) );
  AOI21 U1215 ( .IN1(n593), .IN2(n855), .IN3(n592), .OUT(n594) );
  OAI21 U1216 ( .IN1(n658), .IN2(n688), .IN3(n594), .OUT(n595) );
  AOI21 U1217 ( .IN1(n425), .IN2(n642), .IN3(n595), .OUT(n596) );
  OAI21 U1218 ( .IN1(n905), .IN2(n597), .IN3(n596), .OUT(n598) );
  AOI21 U1219 ( .IN1(n426), .IN2(n599), .IN3(n598), .OUT(n605) );
  AOI22 U1220 ( .IN1(n623), .IN2(n670), .IN3(n669), .IN4(n667), .OUT(n602) );
  AOI22 U1221 ( .IN1(n673), .IN2(n668), .IN3(n680), .IN4(n671), .OUT(n601) );
  AOI22 U1222 ( .IN1(n425), .IN2(n906), .IN3(n603), .IN4(n692), .OUT(n604) );
  OAI21 U1223 ( .IN1(RSTn_BAR), .IN2(n605), .IN3(n604), .OUT(n1064) );
  AOI22 U1224 ( .IN1(n670), .IN2(n426), .IN3(n959), .IN4(n667), .OUT(n607) );
  AOI22 U1225 ( .IN1(n673), .IN2(n958), .IN3(n951), .IN4(n680), .OUT(n606) );
  AOI22 U1226 ( .IN1(n426), .IN2(n646), .IN3(n428), .IN4(n610), .OUT(n609) );
  AOI22 U1227 ( .IN1(n645), .IN2(n427), .IN3(n419), .IN4(n884), .OUT(n608) );
  AOI22 U1228 ( .IN1(n646), .IN2(n420), .IN3(n422), .IN4(n610), .OUT(n612) );
  AOI22 U1229 ( .IN1(n645), .IN2(n421), .IN3(n423), .IN4(n884), .OUT(n611) );
  AOI21 U1230 ( .IN1(n630), .IN2(n1519), .IN3(n613), .OUT(n620) );
  OAI21 U1231 ( .IN1(n423), .IN2(n615), .IN3(n614), .OUT(n617) );
  AOI22 U1232 ( .IN1(n1568), .IN2(Adder_dataout[4]), .IN3(n425), .IN4(n889), 
        .OUT(n616) );
  OAI21 U1233 ( .IN1(n893), .IN2(n617), .IN3(n616), .OUT(n618) );
  AOI21 U1234 ( .IN1(n668), .IN2(n897), .IN3(n618), .OUT(n619) );
  OAI21 U1235 ( .IN1(n621), .IN2(n620), .IN3(n619), .OUT(n622) );
  AOI21 U1236 ( .IN1(n679), .IN2(n629), .IN3(n622), .OUT(n628) );
  AOI22 U1237 ( .IN1(n670), .IN2(n686), .IN3(n623), .IN4(n667), .OUT(n625) );
  AOI22 U1238 ( .IN1(n673), .IN2(n669), .IN3(n680), .IN4(n668), .OUT(n624) );
  AOI22 U1239 ( .IN1(n423), .IN2(n694), .IN3(n626), .IN4(n692), .OUT(n627) );
  OAI21 U1240 ( .IN1(RSTn_BAR), .IN2(n628), .IN3(n627), .OUT(n1065) );
  AOI22 U1241 ( .IN1(n1568), .IN2(Adder_dataout[0]), .IN3(n420), .IN4(n889), 
        .OUT(n631) );
  OAI21 U1242 ( .IN1(n419), .IN2(n893), .IN3(n631), .OUT(n632) );
  AOI21 U1243 ( .IN1(n897), .IN2(n951), .IN3(n632), .OUT(n633) );
  OAI21 U1244 ( .IN1(n689), .IN2(n634), .IN3(n633), .OUT(n635) );
  AOI22 U1245 ( .IN1(n419), .IN2(n694), .IN3(n429), .IN4(n635), .OUT(n636) );
  OAI21 U1246 ( .IN1(n637), .IN2(n879), .IN3(n636), .OUT(n1069) );
  NOR2X1 U1247 ( .IN1(n893), .IN2(n891), .OUT(n643) );
  MUX2X1 U1248 ( .IN1(n643), .IN2(n642), .S(n424), .OUT(n661) );
  AOI22 U1249 ( .IN1(n646), .IN2(n422), .IN3(n423), .IN4(n645), .OUT(n647) );
  OAI21 U1250 ( .IN1(n314), .IN2(n648), .IN3(n647), .OUT(n656) );
  AOI22 U1251 ( .IN1(n1568), .IN2(Adder_dataout[6]), .IN3(
        Final_Mantissa_reg[10]), .IN4(n889), .OUT(n654) );
  MUX2X1 U1252 ( .IN1(n427), .IN2(n426), .S(n1482), .OUT(n650) );
  NOR2X1 U1253 ( .IN1(n1519), .IN2(n1498), .OUT(n649) );
  NAND3X1 U1254 ( .IN1(n866), .IN2(n864), .IN3(n865), .OUT(n652) );
  NAND3X1 U1255 ( .IN1(n654), .IN2(n653), .IN3(n652), .OUT(n655) );
  AOI21 U1256 ( .IN1(n855), .IN2(n656), .IN3(n655), .OUT(n657) );
  OAI21 U1257 ( .IN1(n659), .IN2(n658), .IN3(n657), .OUT(n660) );
  NOR2X1 U1258 ( .IN1(n661), .IN2(n660), .OUT(n662) );
  OAI21 U1259 ( .IN1(n905), .IN2(n663), .IN3(n662), .OUT(n665) );
  AOI21 U1260 ( .IN1(n867), .IN2(n666), .IN3(n665), .OUT(n678) );
  AOI22 U1261 ( .IN1(n670), .IN2(n669), .IN3(n668), .IN4(n667), .OUT(n675) );
  AOI22 U1262 ( .IN1(n673), .IN2(n671), .IN3(n680), .IN4(n221), .OUT(n674) );
  AOI22 U1263 ( .IN1(n424), .IN2(n906), .IN3(n676), .IN4(n692), .OUT(n677) );
  OAI21 U1264 ( .IN1(RSTn_BAR), .IN2(n678), .IN3(n677), .OUT(n1063) );
  AOI22 U1265 ( .IN1(n884), .IN2(n681), .IN3(n680), .IN4(n679), .OUT(n682) );
  AOI22 U1266 ( .IN1(n308), .IN2(n420), .IN3(n419), .IN4(n298), .OUT(n684) );
  AOI22 U1267 ( .IN1(n1568), .IN2(Adder_dataout[1]), .IN3(n421), .IN4(n889), 
        .OUT(n683) );
  OAI21 U1268 ( .IN1(n684), .IN2(n893), .IN3(n683), .OUT(n685) );
  AOI21 U1269 ( .IN1(n897), .IN2(n686), .IN3(n685), .OUT(n687) );
  OAI21 U1270 ( .IN1(n689), .IN2(n688), .IN3(n687), .OUT(n690) );
  AOI21 U1271 ( .IN1(n691), .IN2(n426), .IN3(n690), .OUT(n696) );
  AOI22 U1272 ( .IN1(n420), .IN2(n694), .IN3(n693), .IN4(n692), .OUT(n695) );
  OAI21 U1273 ( .IN1(RSTn_BAR), .IN2(n696), .IN3(n695), .OUT(n1068) );
  NANDX2 U1274 ( .IN1(n429), .IN2(n1569), .OUT(n1625) );
  NOR2X1 U1275 ( .IN1(n301), .IN2(n1580), .OUT(n1567) );
  OAI21 U1276 ( .IN1(n415), .IN2(n1565), .IN3(n429), .OUT(n1260) );
  NOR2X1 U1277 ( .IN1(StateMC[2]), .IN2(n1626), .OUT(n699) );
  OAI21 U1278 ( .IN1(n1556), .IN2(n700), .IN3(n699), .OUT(n701) );
  OAI21 U1279 ( .IN1(n1568), .IN2(n701), .IN3(n429), .OUT(n702) );
  NOR2X1 U1280 ( .IN1(n1548), .IN2(n1625), .OUT(n1562) );
  OAI21 U1281 ( .IN1(n802), .IN2(n1562), .IN3(n188), .OUT(n760) );
  OAI21 U1282 ( .IN1(n1321), .IN2(n714), .IN3(N155), .OUT(n704) );
  AOI21 U1283 ( .IN1(n417), .IN2(n716), .IN3(n704), .OUT(n710) );
  NOR2X1 U1284 ( .IN1(N164), .IN2(N165), .OUT(n713) );
  AOI22 U1285 ( .IN1(n713), .IN2(Datain1[1]), .IN3(n225), .IN4(n712), .OUT(
        n709) );
  AOI22 U1286 ( .IN1(n713), .IN2(Datain1[0]), .IN3(n418), .IN4(n712), .OUT(
        n708) );
  OAI21 U1287 ( .IN1(n1312), .IN2(n714), .IN3(DP_OP_982J1_125_6202_n8), .OUT(
        n706) );
  AOI21 U1288 ( .IN1(n716), .IN2(n416), .IN3(n706), .OUT(n707) );
  AOI22 U1289 ( .IN1(n710), .IN2(n709), .IN3(n708), .IN4(n707), .OUT(n726) );
  OAI21 U1290 ( .IN1(DP_OP_982J1_125_6202_n137), .IN2(n714), .IN3(N155), .OUT(
        n711) );
  AOI21 U1291 ( .IN1(Datain1[13]), .IN2(n716), .IN3(n711), .OUT(n720) );
  AOI22 U1292 ( .IN1(n713), .IN2(Datain1[9]), .IN3(Datain1[15]), .IN4(n712), 
        .OUT(n719) );
  AOI22 U1293 ( .IN1(n713), .IN2(Datain1[8]), .IN3(Datain1[14]), .IN4(n712), 
        .OUT(n718) );
  OAI21 U1294 ( .IN1(n259), .IN2(n714), .IN3(DP_OP_982J1_125_6202_n8), .OUT(
        n715) );
  AOI21 U1295 ( .IN1(Datain1[12]), .IN2(n716), .IN3(n715), .OUT(n717) );
  AOI22 U1296 ( .IN1(n720), .IN2(n719), .IN3(n718), .IN4(n717), .OUT(n721) );
  INVX4 U1297 ( .IN(N419), .OUT(n1411) );
  INVX4 U1298 ( .IN(N420), .OUT(n1345) );
  NOR2X1 U1299 ( .IN1(N424), .IN2(N425), .OUT(n722) );
  AOI21 U1300 ( .IN1(n724), .IN2(N166), .IN3(n723), .OUT(n725) );
  OAI21 U1301 ( .IN1(N166), .IN2(n726), .IN3(n725), .OUT(n759) );
  OAI21 U1302 ( .IN1(n827), .IN2(n740), .IN3(N151), .OUT(n730) );
  AOI21 U1303 ( .IN1(Datain2[5]), .IN2(n742), .IN3(n730), .OUT(n736) );
  NOR2X1 U1304 ( .IN1(N152), .IN2(N153), .OUT(n739) );
  AOI22 U1305 ( .IN1(n739), .IN2(Datain2[1]), .IN3(Datain2[7]), .IN4(n738), 
        .OUT(n735) );
  AOI22 U1306 ( .IN1(n739), .IN2(Datain2[0]), .IN3(Datain2[6]), .IN4(n738), 
        .OUT(n734) );
  OAI21 U1307 ( .IN1(n830), .IN2(n740), .IN3(DP_OP_981J1_124_6202_n8), .OUT(
        n732) );
  AOI21 U1308 ( .IN1(n742), .IN2(Datain2[4]), .IN3(n732), .OUT(n733) );
  AOI22 U1309 ( .IN1(n736), .IN2(n735), .IN3(n734), .IN4(n733), .OUT(n757) );
  OAI21 U1310 ( .IN1(DP_OP_981J1_124_6202_n137), .IN2(n740), .IN3(N151), .OUT(
        n737) );
  AOI21 U1311 ( .IN1(DP_OP_982J1_125_6202_n181), .IN2(n742), .IN3(n737), .OUT(
        n746) );
  AOI22 U1312 ( .IN1(n739), .IN2(DP_OP_982J1_125_6202_n177), .IN3(Datain2[15]), 
        .IN4(n738), .OUT(n745) );
  AOI22 U1313 ( .IN1(n739), .IN2(Datain2[8]), .IN3(DP_OP_982J1_125_6202_n182), 
        .IN4(n738), .OUT(n744) );
  OAI21 U1314 ( .IN1(n1570), .IN2(n740), .IN3(DP_OP_981J1_124_6202_n8), .OUT(
        n741) );
  AOI21 U1315 ( .IN1(DP_OP_982J1_125_6202_n180), .IN2(n742), .IN3(n741), .OUT(
        n743) );
  AOI22 U1316 ( .IN1(n746), .IN2(n745), .IN3(n744), .IN4(n743), .OUT(n747) );
  NOR2X1 U1317 ( .IN1(N366), .IN2(N365), .OUT(n749) );
  NOR2X1 U1318 ( .IN1(N368), .IN2(N369), .OUT(n750) );
  AOI22 U1319 ( .IN1(n1357), .IN2(N363), .IN3(n197), .IN4(n772), .OUT(n754) );
  AOI21 U1320 ( .IN1(n755), .IN2(N154), .IN3(n754), .OUT(n756) );
  OAI21 U1321 ( .IN1(N154), .IN2(n757), .IN3(n756), .OUT(n758) );
  NAND3X1 U1322 ( .IN1(n760), .IN2(n759), .IN3(n758), .OUT(n1071) );
  AOI22 U1323 ( .IN1(n861), .IN2(add_x_35_A_0_), .IN3(add_x_35_A_1_), .IN4(
        n188), .OUT(n761) );
  AOI22 U1324 ( .IN1(n802), .IN2(n861), .IN3(n762), .IN4(n1562), .OUT(n800) );
  OAI21 U1325 ( .IN1(n827), .IN2(n770), .IN3(N147), .OUT(n764) );
  NOR2X1 U1326 ( .IN1(N148), .IN2(N149), .OUT(n768) );
  OAI21 U1327 ( .IN1(n830), .IN2(n770), .IN3(n769), .OUT(n766) );
  INVX4 U1328 ( .IN(N363), .OUT(n1397) );
  INVX4 U1329 ( .IN(n772), .OUT(n1443) );
  OAI21 U1330 ( .IN1(n1321), .IN2(n786), .IN3(n202), .OUT(n776) );
  AOI21 U1331 ( .IN1(n417), .IN2(n788), .IN3(n776), .OUT(n782) );
  NOR2X1 U1332 ( .IN1(N160), .IN2(N161), .OUT(n785) );
  AOI22 U1333 ( .IN1(n785), .IN2(Datain1[1]), .IN3(n225), .IN4(n784), .OUT(
        n781) );
  AOI22 U1334 ( .IN1(n785), .IN2(Datain1[0]), .IN3(n418), .IN4(n784), .OUT(
        n780) );
  OAI21 U1335 ( .IN1(n1312), .IN2(n786), .IN3(n198), .OUT(n778) );
  AOI21 U1336 ( .IN1(n416), .IN2(n788), .IN3(n778), .OUT(n779) );
  AOI22 U1337 ( .IN1(n782), .IN2(n781), .IN3(n780), .IN4(n779), .OUT(n798) );
  OAI21 U1338 ( .IN1(DP_OP_982J1_125_6202_n137), .IN2(n786), .IN3(n202), .OUT(
        n783) );
  AOI21 U1339 ( .IN1(Datain1[13]), .IN2(n788), .IN3(n783), .OUT(n792) );
  AOI22 U1340 ( .IN1(n785), .IN2(Datain1[9]), .IN3(Datain1[15]), .IN4(n784), 
        .OUT(n791) );
  AOI22 U1341 ( .IN1(n785), .IN2(Datain1[8]), .IN3(Datain1[14]), .IN4(n784), 
        .OUT(n790) );
  OAI21 U1342 ( .IN1(n259), .IN2(n786), .IN3(n198), .OUT(n787) );
  AOI21 U1343 ( .IN1(Datain1[12]), .IN2(n788), .IN3(n787), .OUT(n789) );
  AOI22 U1344 ( .IN1(n792), .IN2(n791), .IN3(n790), .IN4(n789), .OUT(n793) );
  OAI21 U1345 ( .IN1(n1323), .IN2(n794), .IN3(n1564), .OUT(n795) );
  AOI21 U1346 ( .IN1(n796), .IN2(N162), .IN3(n795), .OUT(n797) );
  OAI21 U1347 ( .IN1(N162), .IN2(n798), .IN3(n797), .OUT(n799) );
  NOR2X1 U1348 ( .IN1(n189), .IN2(n1479), .OUT(n1475) );
  AOI21 U1349 ( .IN1(n189), .IN2(n1479), .IN3(n1475), .OUT(n801) );
  AOI22 U1350 ( .IN1(n802), .IN2(n189), .IN3(n801), .IN4(n1562), .OUT(n852) );
  OAI21 U1351 ( .IN1(n1321), .IN2(n814), .IN3(N155), .OUT(n804) );
  AOI21 U1352 ( .IN1(n417), .IN2(n816), .IN3(n804), .OUT(n810) );
  NOR2X1 U1353 ( .IN1(N156), .IN2(N157), .OUT(n813) );
  AOI22 U1354 ( .IN1(n813), .IN2(Datain1[1]), .IN3(n225), .IN4(n812), .OUT(
        n809) );
  AOI22 U1355 ( .IN1(Datain1[0]), .IN2(n813), .IN3(n418), .IN4(n812), .OUT(
        n808) );
  OAI21 U1356 ( .IN1(n1312), .IN2(n814), .IN3(DP_OP_982J1_125_6202_n8), .OUT(
        n806) );
  AOI21 U1357 ( .IN1(n416), .IN2(n816), .IN3(n806), .OUT(n807) );
  AOI22 U1358 ( .IN1(n810), .IN2(n809), .IN3(n808), .IN4(n807), .OUT(n824) );
  OAI21 U1359 ( .IN1(DP_OP_982J1_125_6202_n137), .IN2(n814), .IN3(N155), .OUT(
        n811) );
  AOI21 U1360 ( .IN1(Datain1[13]), .IN2(n816), .IN3(n811), .OUT(n820) );
  AOI22 U1361 ( .IN1(Datain1[9]), .IN2(n813), .IN3(Datain1[15]), .IN4(n812), 
        .OUT(n819) );
  AOI22 U1362 ( .IN1(n813), .IN2(Datain1[8]), .IN3(Datain1[14]), .IN4(n812), 
        .OUT(n818) );
  OAI21 U1363 ( .IN1(n259), .IN2(n814), .IN3(DP_OP_982J1_125_6202_n8), .OUT(
        n815) );
  AOI21 U1364 ( .IN1(Datain1[12]), .IN2(n816), .IN3(n815), .OUT(n817) );
  AOI22 U1365 ( .IN1(n820), .IN2(n819), .IN3(n818), .IN4(n817), .OUT(n821) );
  AOI21 U1366 ( .IN1(n822), .IN2(N158), .IN3(n1318), .OUT(n823) );
  OAI21 U1367 ( .IN1(N158), .IN2(n824), .IN3(n823), .OUT(n851) );
  OAI21 U1368 ( .IN1(n827), .IN2(n839), .IN3(N151), .OUT(n828) );
  AOI21 U1369 ( .IN1(Datain2[5]), .IN2(n841), .IN3(n828), .OUT(n835) );
  NOR2X1 U1370 ( .IN1(N144), .IN2(N145), .OUT(n838) );
  AOI22 U1371 ( .IN1(n838), .IN2(Datain2[1]), .IN3(Datain2[7]), .IN4(n837), 
        .OUT(n834) );
  AOI22 U1372 ( .IN1(n838), .IN2(Datain2[0]), .IN3(Datain2[6]), .IN4(n837), 
        .OUT(n833) );
  OAI21 U1373 ( .IN1(n830), .IN2(n839), .IN3(DP_OP_981J1_124_6202_n8), .OUT(
        n831) );
  AOI21 U1374 ( .IN1(Datain2[4]), .IN2(n841), .IN3(n831), .OUT(n832) );
  AOI22 U1375 ( .IN1(n835), .IN2(n834), .IN3(n833), .IN4(n832), .OUT(n847) );
  OAI21 U1376 ( .IN1(DP_OP_981J1_124_6202_n137), .IN2(n839), .IN3(N151), .OUT(
        n836) );
  AOI21 U1377 ( .IN1(DP_OP_982J1_125_6202_n181), .IN2(n841), .IN3(n836), .OUT(
        n845) );
  AOI22 U1378 ( .IN1(n838), .IN2(DP_OP_982J1_125_6202_n177), .IN3(Datain2[15]), 
        .IN4(n837), .OUT(n844) );
  AOI22 U1379 ( .IN1(Datain2[8]), .IN2(n838), .IN3(DP_OP_982J1_125_6202_n182), 
        .IN4(n837), .OUT(n843) );
  OAI21 U1380 ( .IN1(n1570), .IN2(n839), .IN3(DP_OP_981J1_124_6202_n8), .OUT(
        n840) );
  AOI21 U1381 ( .IN1(DP_OP_982J1_125_6202_n180), .IN2(n841), .IN3(n840), .OUT(
        n842) );
  AOI22 U1382 ( .IN1(n845), .IN2(n844), .IN3(n843), .IN4(n842), .OUT(n846) );
  MUX2X1 U1383 ( .IN1(n847), .IN2(n846), .S(N146), .OUT(n848) );
  OAI21 U1384 ( .IN1(n1357), .IN2(n849), .IN3(n848), .OUT(n850) );
  NAND3X1 U1385 ( .IN1(n852), .IN2(n851), .IN3(n850), .OUT(n1072) );
  AOI22 U1386 ( .IN1(n1568), .IN2(n189), .IN3(n419), .IN4(n889), .OUT(n853) );
  OAI21 U1387 ( .IN1(n1298), .IN2(n312), .IN3(n853), .OUT(n854) );
  AOI21 U1388 ( .IN1(n897), .IN2(n958), .IN3(n854), .OUT(n859) );
  NAND3X1 U1389 ( .IN1(n859), .IN2(n858), .IN3(n857), .OUT(n860) );
  AOI22 U1390 ( .IN1(n428), .IN2(n876), .IN3(n429), .IN4(n860), .OUT(n664) );
  AOI22 U1391 ( .IN1(n1568), .IN2(n861), .IN3(n428), .IN4(n889), .OUT(n862) );
  OAI21 U1392 ( .IN1(n1298), .IN2(n299), .IN3(n862), .OUT(n863) );
  AOI21 U1393 ( .IN1(n897), .IN2(n959), .IN3(n863), .OUT(n871) );
  NAND3X1 U1394 ( .IN1(n866), .IN2(n1531), .IN3(n865), .OUT(n870) );
  NAND3X1 U1395 ( .IN1(n871), .IN2(n870), .IN3(n869), .OUT(n872) );
  AOI22 U1396 ( .IN1(n427), .IN2(n876), .IN3(n429), .IN4(n872), .OUT(n672) );
  NOR2X1 U1397 ( .IN1(RSTn_BAR), .IN2(n299), .OUT(n873) );
  AOI22 U1398 ( .IN1(n913), .IN2(n188), .IN3(n873), .IN4(n889), .OUT(n883) );
  NAND3X1 U1399 ( .IN1(n1298), .IN2(n875), .IN3(n874), .OUT(n877) );
  AOI21 U1400 ( .IN1(n877), .IN2(n429), .IN3(n876), .OUT(n878) );
  OAI21 U1401 ( .IN1(n880), .IN2(n879), .IN3(n878), .OUT(n881) );
  NAND3X1 U1402 ( .IN1(n885), .IN2(n296), .IN3(n884), .OUT(n887) );
  OAI21 U1403 ( .IN1(n887), .IN2(n886), .IN3(n1499), .OUT(n888) );
  NAND3X1 U1404 ( .IN1(n1223), .IN2(n888), .IN3(n1530), .OUT(n902) );
  AOI22 U1405 ( .IN1(n1568), .IN2(Adder_dataout[7]), .IN3(carry_reg), .IN4(
        n889), .OUT(n900) );
  OAI21 U1406 ( .IN1(n310), .IN2(n891), .IN3(n296), .OUT(n895) );
  NOR2X1 U1407 ( .IN1(n892), .IN2(n891), .OUT(n907) );
  NOR2X1 U1408 ( .IN1(n893), .IN2(n907), .OUT(n894) );
  AOI22 U1409 ( .IN1(n897), .IN2(n896), .IN3(n895), .IN4(n894), .OUT(n898) );
  NAND3X1 U1410 ( .IN1(n1627), .IN2(n911), .IN3(n910), .OUT(n912) );
  AOI22 U1411 ( .IN1(n913), .IN2(Adder_carryout), .IN3(carry_reg), .IN4(n912), 
        .OUT(n914) );
  OAI21 U1412 ( .IN1(n1308), .IN2(n1300), .IN3(n914), .OUT(n1061) );
  NOR2X1 U1413 ( .IN1(Final_Exponent_reg[4]), .IN2(Final_Exponent_reg[7]), 
        .OUT(n916) );
  NAND3X1 U1414 ( .IN1(n295), .IN2(n304), .IN3(n916), .OUT(n917) );
  AOI21 U1415 ( .IN1(n1257), .IN2(n1274), .IN3(n1627), .OUT(n925) );
  NOR2X1 U1416 ( .IN1(n925), .IN2(n924), .OUT(n926) );
  INVX4 U1417 ( .IN(n926), .OUT(n1179) );
  AOI22 U1418 ( .IN1(n411), .IN2(n1179), .IN3(DP_OP_982J1_125_6202_n177), 
        .IN4(n1564), .OUT(n1047) );
  OAI21 U1419 ( .IN1(Final_Exponent_reg[1]), .IN2(Final_Exponent_reg[2]), 
        .IN3(DP_OP_979_173_2805_n76), .OUT(n931) );
  AOI22 U1420 ( .IN1(n426), .IN2(n1227), .IN3(n427), .IN4(n1203), .OUT(n933)
         );
  AOI22 U1421 ( .IN1(n1205), .IN2(n992), .IN3(n935), .IN4(n934), .OUT(n939) );
  OAI21 U1422 ( .IN1(n410), .IN2(n942), .IN3(n1003), .OUT(n1234) );
  NOR2X1 U1423 ( .IN1(n1487), .IN2(n1234), .OUT(n1017) );
  OAI21 U1424 ( .IN1(n999), .IN2(n1210), .IN3(n994), .OUT(n943) );
  NAND3X1 U1425 ( .IN1(n951), .IN2(n950), .IN3(n975), .OUT(n956) );
  AOI21 U1426 ( .IN1(n956), .IN2(n955), .IN3(n954), .OUT(n1014) );
  NAND3X1 U1427 ( .IN1(n414), .IN2(n957), .IN3(n1025), .OUT(n969) );
  AOI22 U1428 ( .IN1(n1227), .IN2(n427), .IN3(n992), .IN4(n958), .OUT(n961) );
  NOR2X1 U1429 ( .IN1(n969), .IN2(n968), .OUT(n970) );
  AOI21 U1430 ( .IN1(n1040), .IN2(n971), .IN3(n970), .OUT(n972) );
  OAI21 U1431 ( .IN1(n1041), .IN2(n1037), .IN3(n972), .OUT(n1186) );
  OAI21 U1432 ( .IN1(n1485), .IN2(n1232), .IN3(n973), .OUT(n974) );
  NOR2X1 U1433 ( .IN1(n1235), .IN2(n1233), .OUT(n982) );
  AOI22 U1434 ( .IN1(n984), .IN2(n983), .IN3(n982), .IN4(n981), .OUT(n985) );
  AOI22 U1435 ( .IN1(n1271), .IN2(C1_DATA14_2), .IN3(C1_DATA6_2), .IN4(n1181), 
        .OUT(n986) );
  OAI21 U1436 ( .IN1(n1184), .IN2(n987), .IN3(n986), .OUT(n988) );
  AOI21 U1437 ( .IN1(C1_DATA2_2), .IN2(n1186), .IN3(n988), .OUT(n1035) );
  NAND3X1 U1438 ( .IN1(n995), .IN2(n414), .IN3(n1247), .OUT(n996) );
  AOI22 U1439 ( .IN1(n1188), .IN2(n411), .IN3(C1_DATA3_2), .IN4(n1187), .OUT(
        n1021) );
  OAI21 U1440 ( .IN1(n1500), .IN2(n1013), .IN3(n1001), .OUT(n1002) );
  OAI21 U1441 ( .IN1(n1485), .IN2(n1505), .IN3(n1005), .OUT(n1006) );
  AOI22 U1442 ( .IN1(n1190), .IN2(n293), .IN3(C1_DATA9_2), .IN4(n1189), .OUT(
        n1020) );
  OAI21 U1443 ( .IN1(n1485), .IN2(n1226), .IN3(n1009), .OUT(n1278) );
  NOR2X1 U1444 ( .IN1(n1014), .IN2(n1013), .OUT(n1030) );
  AOI22 U1445 ( .IN1(n1017), .IN2(n1016), .IN3(n1015), .IN4(n1030), .OUT(n1018) );
  AOI22 U1446 ( .IN1(n1192), .IN2(C1_DATA10_2), .IN3(C1_DATA5_2), .IN4(n1191), 
        .OUT(n1019) );
  NAND3X1 U1447 ( .IN1(n1021), .IN2(n1020), .IN3(n1019), .OUT(n1022) );
  OAI21 U1448 ( .IN1(n1027), .IN2(n1246), .IN3(n1026), .OUT(n1028) );
  NOR2X1 U1449 ( .IN1(n1029), .IN2(n1028), .OUT(n1031) );
  NAND3X1 U1450 ( .IN1(n1035), .IN2(n1034), .IN3(n1033), .OUT(n1036) );
  AOI21 U1451 ( .IN1(n1272), .IN2(C1_DATA12_2), .IN3(n1036), .OUT(n1044) );
  INVX4 U1452 ( .IN(n1039), .OUT(n1199) );
  INVX4 U1453 ( .IN(n1042), .OUT(n1198) );
  AOI22 U1454 ( .IN1(C1_DATA11_2), .IN2(n1199), .IN3(n1198), .IN4(C1_DATA13_2), 
        .OUT(n1043) );
  AOI21 U1455 ( .IN1(n1044), .IN2(n1043), .IN3(n1627), .OUT(n1045) );
  AOI22 U1456 ( .IN1(n1271), .IN2(C1_DATA14_3), .IN3(C1_DATA6_3), .IN4(n1181), 
        .OUT(n1048) );
  OAI21 U1457 ( .IN1(n1184), .IN2(n1049), .IN3(n1048), .OUT(n1050) );
  AOI21 U1458 ( .IN1(C1_DATA2_3), .IN2(n1186), .IN3(n1050), .OUT(n1057) );
  AOI22 U1459 ( .IN1(n1188), .IN2(n409), .IN3(C1_DATA3_3), .IN4(n1187), .OUT(
        n1053) );
  AOI22 U1460 ( .IN1(n1190), .IN2(C1_DATA4_3), .IN3(C1_DATA9_3), .IN4(n1189), 
        .OUT(n1052) );
  AOI22 U1461 ( .IN1(n1192), .IN2(C1_DATA10_3), .IN3(C1_DATA5_3), .IN4(n1191), 
        .OUT(n1051) );
  NAND3X1 U1462 ( .IN1(n1053), .IN2(n1052), .IN3(n1051), .OUT(n1054) );
  NAND3X1 U1463 ( .IN1(n1057), .IN2(n1056), .IN3(n1055), .OUT(n1058) );
  AOI21 U1464 ( .IN1(n1272), .IN2(C1_DATA12_3), .IN3(n1058), .OUT(n1102) );
  AOI22 U1465 ( .IN1(C1_DATA11_3), .IN2(n1199), .IN3(n1198), .IN4(C1_DATA13_3), 
        .OUT(n1059) );
  AOI21 U1466 ( .IN1(n1102), .IN2(n1059), .IN3(n1627), .OUT(n1104) );
  AOI22 U1467 ( .IN1(n410), .IN2(n1179), .IN3(Datain2[7]), .IN4(n1564), .OUT(
        n1120) );
  AOI22 U1468 ( .IN1(n1271), .IN2(n396), .IN3(n410), .IN4(n1181), .OUT(n1105)
         );
  OAI21 U1469 ( .IN1(n1184), .IN2(n410), .IN3(n1105), .OUT(n1106) );
  AOI21 U1470 ( .IN1(n410), .IN2(n1186), .IN3(n1106), .OUT(n1113) );
  AOI22 U1471 ( .IN1(n1188), .IN2(n410), .IN3(n396), .IN4(n1187), .OUT(n1109)
         );
  AOI22 U1472 ( .IN1(n1190), .IN2(n410), .IN3(n396), .IN4(n1189), .OUT(n1108)
         );
  AOI22 U1473 ( .IN1(n1192), .IN2(n410), .IN3(n396), .IN4(n1191), .OUT(n1107)
         );
  NAND3X1 U1474 ( .IN1(n1109), .IN2(n1108), .IN3(n1107), .OUT(n1110) );
  NAND3X1 U1475 ( .IN1(n1113), .IN2(n1112), .IN3(n1111), .OUT(n1114) );
  AOI21 U1476 ( .IN1(n1272), .IN2(C1_DATA12_0), .IN3(n1114), .OUT(n1116) );
  AOI22 U1477 ( .IN1(C1_DATA11_0), .IN2(n1199), .IN3(n1198), .IN4(C1_DATA13_0), 
        .OUT(n1115) );
  AOI21 U1478 ( .IN1(n1116), .IN2(n1115), .IN3(n1627), .OUT(n1117) );
  NAND3X1 U1479 ( .IN1(n1120), .IN2(n1119), .IN3(n1118), .OUT(n1094) );
  AOI22 U1480 ( .IN1(DP_OP_979_173_2805_n78), .IN2(n1179), .IN3(
        DP_OP_982J1_125_6202_n180), .IN4(n1564), .OUT(n1137) );
  AOI22 U1481 ( .IN1(n1271), .IN2(C1_DATA14_5), .IN3(C1_DATA6_5), .IN4(n1181), 
        .OUT(n1121) );
  OAI21 U1482 ( .IN1(n1184), .IN2(n1122), .IN3(n1121), .OUT(n1123) );
  AOI21 U1483 ( .IN1(C1_DATA2_5), .IN2(n1186), .IN3(n1123), .OUT(n1130) );
  AOI22 U1484 ( .IN1(n1188), .IN2(C1_DATA8_5), .IN3(C1_DATA3_5), .IN4(n1187), 
        .OUT(n1126) );
  AOI22 U1485 ( .IN1(n1190), .IN2(C1_DATA4_5), .IN3(C1_DATA9_5), .IN4(n1189), 
        .OUT(n1125) );
  AOI22 U1486 ( .IN1(n1192), .IN2(C1_DATA10_5), .IN3(C1_DATA5_5), .IN4(n1191), 
        .OUT(n1124) );
  NAND3X1 U1487 ( .IN1(n1126), .IN2(n1125), .IN3(n1124), .OUT(n1127) );
  NAND3X1 U1488 ( .IN1(n1128), .IN2(n1129), .IN3(n1130), .OUT(n1131) );
  AOI21 U1489 ( .IN1(n1272), .IN2(C1_DATA12_5), .IN3(n1131), .OUT(n1133) );
  AOI22 U1490 ( .IN1(C1_DATA11_5), .IN2(n1199), .IN3(n1198), .IN4(C1_DATA13_5), 
        .OUT(n1132) );
  AOI21 U1491 ( .IN1(n1133), .IN2(n1132), .IN3(n1627), .OUT(n1134) );
  NAND3X1 U1492 ( .IN1(n1137), .IN2(n1136), .IN3(n1135), .OUT(n1099) );
  AOI22 U1493 ( .IN1(n407), .IN2(n1179), .IN3(Datain2[8]), .IN4(n1564), .OUT(
        n1154) );
  AOI22 U1494 ( .IN1(n1271), .IN2(C1_DATA14_1), .IN3(n406), .IN4(n1181), .OUT(
        n1138) );
  OAI21 U1495 ( .IN1(n1184), .IN2(n1139), .IN3(n1138), .OUT(n1140) );
  AOI21 U1496 ( .IN1(n406), .IN2(n1186), .IN3(n1140), .OUT(n1147) );
  AOI22 U1497 ( .IN1(n1188), .IN2(n407), .IN3(C1_DATA3_1), .IN4(n1187), .OUT(
        n1143) );
  AOI22 U1498 ( .IN1(n1190), .IN2(n407), .IN3(C1_DATA9_1), .IN4(n1189), .OUT(
        n1142) );
  AOI22 U1499 ( .IN1(n1192), .IN2(n406), .IN3(C1_DATA5_1), .IN4(n1191), .OUT(
        n1141) );
  NAND3X1 U1500 ( .IN1(n1145), .IN2(n1146), .IN3(n1147), .OUT(n1148) );
  AOI21 U1501 ( .IN1(n1272), .IN2(C1_DATA12_1), .IN3(n1148), .OUT(n1150) );
  AOI22 U1502 ( .IN1(C1_DATA11_1), .IN2(n1199), .IN3(n1198), .IN4(C1_DATA13_1), 
        .OUT(n1149) );
  AOI21 U1503 ( .IN1(n1150), .IN2(n1149), .IN3(n1627), .OUT(n1151) );
  NAND3X1 U1504 ( .IN1(n1154), .IN2(n1153), .IN3(n1152), .OUT(n1095) );
  AOI22 U1505 ( .IN1(DP_OP_979_173_2805_n79), .IN2(n1179), .IN3(
        DP_OP_982J1_125_6202_n181), .IN4(n1564), .OUT(n1165) );
  AOI22 U1506 ( .IN1(n1188), .IN2(C1_DATA8_6), .IN3(C1_DATA3_6), .IN4(n1187), 
        .OUT(n1158) );
  AOI22 U1507 ( .IN1(n1190), .IN2(C1_DATA4_6), .IN3(C1_DATA9_6), .IN4(n1189), 
        .OUT(n1157) );
  AOI22 U1508 ( .IN1(n1192), .IN2(C1_DATA10_6), .IN3(C1_DATA5_6), .IN4(n1191), 
        .OUT(n1156) );
  NAND3X1 U1509 ( .IN1(n1158), .IN2(n1157), .IN3(n1156), .OUT(n1159) );
  AOI22 U1510 ( .IN1(DP_OP_979_173_2805_n77), .IN2(n1179), .IN3(Datain2[11]), 
        .IN4(n1564), .OUT(n1178) );
  AOI22 U1511 ( .IN1(n1271), .IN2(C1_DATA14_4), .IN3(C1_DATA6_4), .IN4(n1181), 
        .OUT(n1166) );
  OAI21 U1512 ( .IN1(n1184), .IN2(n1167), .IN3(n1166), .OUT(n1168) );
  NAND3X1 U1513 ( .IN1(n1171), .IN2(n1170), .IN3(n1169), .OUT(n1172) );
  AOI22 U1514 ( .IN1(C1_DATA11_4), .IN2(n1199), .IN3(n1198), .IN4(C1_DATA13_4), 
        .OUT(n1174) );
  NAND3X1 U1515 ( .IN1(n1178), .IN2(n1177), .IN3(n1176), .OUT(n1098) );
  AOI22 U1516 ( .IN1(DP_OP_979_173_2805_n80), .IN2(n1179), .IN3(
        DP_OP_982J1_125_6202_n182), .IN4(n1564), .OUT(n1180) );
  OAI21 U1517 ( .IN1(n1615), .IN2(n1388), .IN3(n1180), .OUT(n1200) );
  AOI22 U1518 ( .IN1(n1271), .IN2(C1_DATA14_7), .IN3(C1_DATA6_7), .IN4(n1181), 
        .OUT(n1182) );
  OAI21 U1519 ( .IN1(n1184), .IN2(n1183), .IN3(n1182), .OUT(n1185) );
  AOI22 U1520 ( .IN1(n1188), .IN2(C1_DATA8_7), .IN3(C1_DATA3_7), .IN4(n1187), 
        .OUT(n1195) );
  AOI22 U1521 ( .IN1(n1190), .IN2(C1_DATA4_7), .IN3(C1_DATA9_7), .IN4(n1189), 
        .OUT(n1194) );
  AOI22 U1522 ( .IN1(n1192), .IN2(C1_DATA10_7), .IN3(C1_DATA5_7), .IN4(n1191), 
        .OUT(n1193) );
  NAND3X1 U1523 ( .IN1(n1195), .IN2(n1194), .IN3(n1193), .OUT(n1196) );
  AOI21 U1524 ( .IN1(n1201), .IN2(n1279), .IN3(n1532), .OUT(n1209) );
  AOI22 U1525 ( .IN1(n1230), .IN2(n1205), .IN3(n1229), .IN4(n1204), .OUT(n1206) );
  OAI21 U1526 ( .IN1(n1212), .IN2(n1211), .IN3(n1210), .OUT(n1213) );
  AOI21 U1527 ( .IN1(n1214), .IN2(n1246), .IN3(n1213), .OUT(n1222) );
  AOI22 U1528 ( .IN1(n1234), .IN2(n1217), .IN3(n1216), .IN4(n1215), .OUT(n1218) );
  OAI21 U1529 ( .IN1(n1237), .IN2(n1219), .IN3(n1218), .OUT(n1220) );
  AOI21 U1530 ( .IN1(n1223), .IN2(n1266), .IN3(n1276), .OUT(n1224) );
  NOR2X1 U1531 ( .IN1(n1483), .IN2(n1224), .OUT(n1225) );
  OAI21 U1532 ( .IN1(n1227), .IN2(n1226), .IN3(n414), .OUT(n1255) );
  AOI22 U1533 ( .IN1(n1231), .IN2(n1230), .IN3(n1229), .IN4(n1228), .OUT(n1254) );
  AOI22 U1534 ( .IN1(n1236), .IN2(n1235), .IN3(n1503), .IN4(n1234), .OUT(n1249) );
  AOI22 U1535 ( .IN1(n1241), .IN2(n1240), .IN3(n1239), .IN4(n1238), .OUT(n1242) );
  OAI21 U1536 ( .IN1(n1244), .IN2(n1243), .IN3(n1242), .OUT(n1245) );
  AOI21 U1537 ( .IN1(n1247), .IN2(n1246), .IN3(n1245), .OUT(n1248) );
  AOI21 U1538 ( .IN1(n1252), .IN2(n1251), .IN3(n1250), .OUT(n1253) );
  NOR2X1 U1539 ( .IN1(n1255), .IN2(n1284), .OUT(n1267) );
  NOR2X1 U1540 ( .IN1(n1256), .IN2(n1267), .OUT(n1258) );
  OAI21 U1541 ( .IN1(n223), .IN2(n1258), .IN3(n1257), .OUT(n1292) );
  NOR2X1 U1542 ( .IN1(n1259), .IN2(n1260), .OUT(n1286) );
  AOI21 U1543 ( .IN1(StateMC[2]), .IN2(n301), .IN3(RSTn_BAR), .OUT(n1261) );
  NOR2X1 U1544 ( .IN1(Exc_Ack), .IN2(n1260), .OUT(N270) );
  AOI21 U1545 ( .IN1(n1261), .IN2(n1580), .IN3(N270), .OUT(n1262) );
  AOI22 U1546 ( .IN1(Exc_value[1]), .IN2(n1286), .IN3(n320), .IN4(n1285), 
        .OUT(n1263) );
  OAI21 U1547 ( .IN1(n1627), .IN2(n1294), .IN3(n1263), .OUT(n1093) );
  NOR2X1 U1548 ( .IN1(n1264), .IN2(n1271), .OUT(n1265) );
  OAI21 U1549 ( .IN1(n1266), .IN2(n1276), .IN3(n1265), .OUT(n1268) );
  NOR2X1 U1550 ( .IN1(n1268), .IN2(n1267), .OUT(n1269) );
  NOR2X1 U1551 ( .IN1(n222), .IN2(n1269), .OUT(n1295) );
  AOI22 U1552 ( .IN1(Exc_value[2]), .IN2(n1286), .IN3(n302), .IN4(n1285), 
        .OUT(n1270) );
  OAI21 U1553 ( .IN1(n1627), .IN2(n1293), .IN3(n1270), .OUT(n1101) );
  NOR2X1 U1554 ( .IN1(n1272), .IN2(n1271), .OUT(n1273) );
  NAND3X1 U1555 ( .IN1(n1274), .IN2(n1485), .IN3(n1273), .OUT(n1275) );
  OAI21 U1556 ( .IN1(n1499), .IN2(n1275), .IN3(exc_reg_0_), .OUT(n1282) );
  OAI21 U1557 ( .IN1(n1277), .IN2(n1276), .IN3(n1499), .OUT(n1281) );
  NAND3X1 U1558 ( .IN1(n1282), .IN2(n1281), .IN3(n1280), .OUT(n1283) );
  AOI21 U1559 ( .IN1(n1284), .IN2(n414), .IN3(n1283), .OUT(n1291) );
  AOI22 U1560 ( .IN1(n1286), .IN2(Exc_value[0]), .IN3(exc_reg_0_), .IN4(n1285), 
        .OUT(n1287) );
  OAI21 U1561 ( .IN1(n1627), .IN2(n1291), .IN3(n1287), .OUT(n1092) );
  NAND3X1 U1562 ( .IN1(n223), .IN2(n222), .IN3(n317), .OUT(n1289) );
  NAND3X1 U1563 ( .IN1(exc_reg_0_), .IN2(n302), .IN3(n320), .OUT(n1288) );
  OAI21 U1564 ( .IN1(n1538), .IN2(n1290), .IN3(n1577), .OUT(n1584) );
  NAND3X1 U1565 ( .IN1(n1298), .IN2(n1297), .IN3(n1296), .OUT(n1299) );
  AOI21 U1566 ( .IN1(n1563), .IN2(n1300), .IN3(n1299), .OUT(n1301) );
  OAI21 U1567 ( .IN1(n1581), .IN2(n1302), .IN3(n1301), .OUT(n1303) );
  AOI21 U1568 ( .IN1(n1307), .IN2(Op1_Sign_reg), .IN3(n1517), .OUT(n1624) );
  NOR2X1 U1569 ( .IN1(n1310), .IN2(n1581), .OUT(n1311) );
  AOI22 U1570 ( .IN1(n1535), .IN2(n324), .IN3(n1311), .IN4(n414), .OUT(n1623)
         );
  INVX4 U1571 ( .IN(n1316), .OUT(n1406) );
  NOR2X1 U1572 ( .IN1(n1312), .IN2(n1350), .OUT(n1313) );
  MUX2X1 U1573 ( .IN1(Datain2[1]), .IN2(Datain2[3]), .S(N363), .OUT(n1363) );
  AOI22 U1574 ( .IN1(n1446), .IN2(n1313), .IN3(n1351), .IN4(n1363), .OUT(n1343) );
  MUX2X1 U1575 ( .IN1(Datain2[0]), .IN2(Datain2[2]), .S(N363), .OUT(n1339) );
  AOI22 U1576 ( .IN1(n417), .IN2(n202), .IN3(n1457), .IN4(N419), .OUT(n1315)
         );
  NOR2X1 U1577 ( .IN1(n202), .IN2(N419), .OUT(n1378) );
  NOR2X1 U1578 ( .IN1(n1345), .IN2(n1316), .OUT(n1317) );
  AOI22 U1579 ( .IN1(n1465), .IN2(n1477), .IN3(n1436), .IN4(n1386), .OUT(n1337) );
  NOR2X1 U1580 ( .IN1(n1621), .IN2(n1318), .OUT(n1319) );
  MUX2X1 U1581 ( .IN1(Datain1[0]), .IN2(Datain1[2]), .S(N419), .OUT(n1328) );
  MUX2X1 U1582 ( .IN1(n1322), .IN2(n1321), .S(N419), .OUT(n1358) );
  AOI22 U1583 ( .IN1(n418), .IN2(n1377), .IN3(n417), .IN4(n1427), .OUT(n1324)
         );
  MUX2X1 U1584 ( .IN1(n1326), .IN2(n1435), .S(N420), .OUT(n1327) );
  OAI21 U1585 ( .IN1(n1369), .IN2(n1328), .IN3(n1327), .OUT(n1329) );
  MUX2X1 U1586 ( .IN1(n1330), .IN2(n1352), .S(N363), .OUT(n1422) );
  MUX2X1 U1587 ( .IN1(n1422), .IN2(n1353), .S(N362), .OUT(n1334) );
  NOR2X1 U1588 ( .IN1(n1331), .IN2(Datain2[10]), .OUT(n1332) );
  NAND3X1 U1589 ( .IN1(N363), .IN2(n1454), .IN3(n1396), .OUT(n1333) );
  OAI21 U1590 ( .IN1(n1334), .IN2(n1388), .IN3(n1333), .OUT(n1434) );
  AOI22 U1591 ( .IN1(n1384), .IN2(n1335), .IN3(n1389), .IN4(n1434), .OUT(n1336) );
  AOI21 U1592 ( .IN1(n412), .IN2(n1339), .IN3(n1338), .OUT(n1342) );
  NAND3X1 U1593 ( .IN1(n1343), .IN2(n1342), .IN3(n1341), .OUT(n1080) );
  AOI22 U1594 ( .IN1(n415), .IN2(n1477), .IN3(n419), .IN4(n1565), .OUT(n1344)
         );
  MUX2X1 U1595 ( .IN1(Datain1[2]), .IN2(n416), .S(N419), .OUT(n1370) );
  NAND3X1 U1596 ( .IN1(N420), .IN2(n1444), .IN3(n1384), .OUT(n1346) );
  OAI21 U1597 ( .IN1(n1347), .IN2(n1426), .IN3(n1346), .OUT(n1368) );
  NAND3X1 U1598 ( .IN1(n1350), .IN2(n1349), .IN3(n1348), .OUT(n1445) );
  AOI22 U1599 ( .IN1(n1465), .IN2(n1552), .IN3(n1445), .IN4(n1386), .OUT(n1366) );
  MUX2X1 U1600 ( .IN1(Datain2[2]), .IN2(Datain2[4]), .S(N363), .OUT(n1395) );
  NOR2X1 U1601 ( .IN1(n1352), .IN2(N363), .OUT(n1390) );
  OAI21 U1602 ( .IN1(n1397), .IN2(n1462), .IN3(n1355), .OUT(n1356) );
  AOI22 U1603 ( .IN1(n1357), .IN2(n1390), .IN3(n769), .IN4(n1356), .OUT(n1441)
         );
  NAND3X1 U1604 ( .IN1(n1379), .IN2(n1359), .IN3(n1384), .OUT(n1360) );
  OAI21 U1605 ( .IN1(n1441), .IN2(n1361), .IN3(n1360), .OUT(n1362) );
  AOI21 U1606 ( .IN1(n412), .IN2(n1363), .IN3(n1362), .OUT(n1364) );
  NAND3X1 U1607 ( .IN1(n1366), .IN2(n1365), .IN3(n1364), .OUT(n1367) );
  AOI21 U1608 ( .IN1(n1369), .IN2(n1368), .IN3(n1367), .OUT(n1373) );
  MUX2X1 U1609 ( .IN1(n1371), .IN2(n1412), .S(n202), .OUT(n1372) );
  AOI22 U1610 ( .IN1(n415), .IN2(n1552), .IN3(n420), .IN4(n1565), .OUT(n1374)
         );
  MUX2X1 U1611 ( .IN1(Datain1[3]), .IN2(n417), .S(N419), .OUT(n1417) );
  AOI22 U1612 ( .IN1(n1377), .IN2(n1376), .IN3(n202), .IN4(n1375), .OUT(n1382)
         );
  NOR2X1 U1613 ( .IN1(Datain1[2]), .IN2(N419), .OUT(n1380) );
  AOI22 U1614 ( .IN1(N420), .IN2(n1450), .IN3(n1380), .IN4(n1379), .OUT(n1381)
         );
  AOI22 U1615 ( .IN1(n1465), .IN2(n1554), .IN3(n1385), .IN4(n1384), .OUT(n1393) );
  NAND3X1 U1616 ( .IN1(n418), .IN2(n1411), .IN3(n1386), .OUT(n1392) );
  AOI21 U1617 ( .IN1(N362), .IN2(n355), .IN3(n1388), .OUT(n1455) );
  NAND3X1 U1618 ( .IN1(n1390), .IN2(n1455), .IN3(n1389), .OUT(n1391) );
  NAND3X1 U1619 ( .IN1(n1393), .IN2(n1392), .IN3(n1391), .OUT(n1394) );
  AOI21 U1620 ( .IN1(n412), .IN2(n1395), .IN3(n1394), .OUT(n1415) );
  NAND3X1 U1621 ( .IN1(Datain2[5]), .IN2(N363), .IN3(n197), .OUT(n1399) );
  AOI22 U1622 ( .IN1(n1402), .IN2(n1401), .IN3(n1400), .IN4(n1443), .OUT(n1403) );
  OAI21 U1623 ( .IN1(n1404), .IN2(n1453), .IN3(n1403), .OUT(n1424) );
  NAND3X1 U1624 ( .IN1(Datain1[3]), .IN2(n1406), .IN3(n1405), .OUT(n1407) );
  AOI22 U1625 ( .IN1(n1411), .IN2(n1410), .IN3(n417), .IN4(n1409), .OUT(n1430)
         );
  MUX2X1 U1626 ( .IN1(n1430), .IN2(n1412), .S(n198), .OUT(n1413) );
  NAND3X1 U1627 ( .IN1(n1415), .IN2(n1414), .IN3(n1413), .OUT(n1078) );
  AOI22 U1628 ( .IN1(n415), .IN2(n1554), .IN3(n421), .IN4(n1565), .OUT(n1416)
         );
  AOI22 U1629 ( .IN1(n198), .IN2(n1417), .IN3(n416), .IN4(n1427), .OUT(n1418)
         );
  AOI22 U1630 ( .IN1(n315), .IN2(n1465), .IN3(n1419), .IN4(n1451), .OUT(n1420)
         );
  OAI21 U1631 ( .IN1(n1422), .IN2(n1421), .IN3(n1420), .OUT(n1423) );
  AOI21 U1632 ( .IN1(n769), .IN2(n1424), .IN3(n1423), .OUT(n1432) );
  OAI21 U1633 ( .IN1(n1427), .IN2(n1426), .IN3(n1425), .OUT(n1428) );
  AOI22 U1634 ( .IN1(n1456), .IN2(n416), .IN3(n418), .IN4(n1428), .OUT(n1429)
         );
  MUX2X1 U1635 ( .IN1(n1430), .IN2(n1429), .S(n202), .OUT(n1431) );
  AOI22 U1636 ( .IN1(n415), .IN2(n315), .IN3(n422), .IN4(n1565), .OUT(n1433)
         );
  AOI22 U1637 ( .IN1(n1465), .IN2(n316), .IN3(n1434), .IN4(n1443), .OUT(n1439)
         );
  NAND3X1 U1638 ( .IN1(n1439), .IN2(n1438), .IN3(n1437), .OUT(n1076) );
  AOI22 U1639 ( .IN1(n415), .IN2(n316), .IN3(n423), .IN4(n1565), .OUT(n1440)
         );
  AOI22 U1640 ( .IN1(n1465), .IN2(n318), .IN3(n1443), .IN4(n1442), .OUT(n1448)
         );
  AOI22 U1641 ( .IN1(n1446), .IN2(n1445), .IN3(n1451), .IN4(n1444), .OUT(n1447) );
  AOI22 U1642 ( .IN1(n415), .IN2(n318), .IN3(n425), .IN4(n1565), .OUT(n1449)
         );
  AOI22 U1643 ( .IN1(n1465), .IN2(n319), .IN3(n1452), .IN4(n1451), .OUT(n1460)
         );
  NAND3X1 U1644 ( .IN1(n1455), .IN2(n1454), .IN3(n1463), .OUT(n1459) );
  NAND3X1 U1645 ( .IN1(n1460), .IN2(n1459), .IN3(n1458), .OUT(n1074) );
  AOI22 U1646 ( .IN1(n415), .IN2(n319), .IN3(n424), .IN4(n1565), .OUT(n1461)
         );
  NOR2X1 U1647 ( .IN1(N362), .IN2(n1462), .OUT(n1464) );
  AOI22 U1648 ( .IN1(Op2_Mantissa_reg_7_), .IN2(n1465), .IN3(n1464), .IN4(
        n1463), .OUT(n1466) );
  OAI21 U1649 ( .IN1(n202), .IN2(n1467), .IN3(n1466), .OUT(n1073) );
  AOI22 U1650 ( .IN1(n415), .IN2(Op2_Mantissa_reg_7_), .IN3(n410), .IN4(n1565), 
        .OUT(ExcCheck_Datain_7__BAR) );
  AOI22 U1651 ( .IN1(n415), .IN2(n410), .IN3(n407), .IN4(n1565), .OUT(n1469)
         );
  AOI22 U1652 ( .IN1(n415), .IN2(n407), .IN3(n411), .IN4(n1565), .OUT(n1470)
         );
  AOI22 U1653 ( .IN1(n415), .IN2(n411), .IN3(DP_OP_979_173_2805_n76), .IN4(
        n1565), .OUT(ExcCheck_Datain_10__BAR) );
  AOI22 U1654 ( .IN1(n415), .IN2(DP_OP_979_173_2805_n76), .IN3(
        DP_OP_979_173_2805_n77), .IN4(n1565), .OUT(n1472) );
  AOI22 U1655 ( .IN1(n415), .IN2(DP_OP_979_173_2805_n77), .IN3(
        DP_OP_979_173_2805_n78), .IN4(n1565), .OUT(n1473) );
  AOI22 U1656 ( .IN1(n415), .IN2(DP_OP_979_173_2805_n78), .IN3(
        DP_OP_979_173_2805_n79), .IN4(n1565), .OUT(ExcCheck_Datain_13__BAR) );
  AOI22 U1657 ( .IN1(n415), .IN2(DP_OP_979_173_2805_n79), .IN3(
        DP_OP_979_173_2805_n80), .IN4(n1565), .OUT(n1474) );
  NOR2X1 U1658 ( .IN1(n1475), .IN2(n1548), .OUT(n1476) );
  MUX2X1 U1659 ( .IN1(add_x_35_A_3_), .IN2(n1477), .S(n1476), .OUT(n1478) );
  NOR2X1 U1660 ( .IN1(n1625), .IN2(n1478), .OUT(n116) );
  MUX2X1 U1661 ( .IN1(n1552), .IN2(add_x_35_A_4_), .S(n1480), .OUT(n1481) );
  NOR2X1 U1662 ( .IN1(n1481), .IN2(n1625), .OUT(n117) );
  OAI21 U1663 ( .IN1(n219), .IN2(n413), .IN3(n1608), .OUT(n1089) );
  NOR2X1 U1664 ( .IN1(n219), .IN2(n1625), .OUT(N252) );
  OAI21 U1665 ( .IN1(n218), .IN2(n413), .IN3(n1609), .OUT(n1088) );
  NOR2X1 U1666 ( .IN1(n218), .IN2(n1625), .OUT(N253) );
  AOI22 U1667 ( .IN1(n1588), .IN2(Debug_reg[0]), .IN3(StateMC[0]), .IN4(n1587), 
        .OUT(n1486) );
  NAND3X1 U1668 ( .IN1(n277), .IN2(n1488), .IN3(n1487), .OUT(n1489) );
  NAND3X1 U1669 ( .IN1(n1492), .IN2(n1491), .IN3(n1490), .OUT(n1496) );
  OAI21 U1670 ( .IN1(n1496), .IN2(n1495), .IN3(n1494), .OUT(n1497) );
  AOI21 U1671 ( .IN1(n1499), .IN2(n1498), .IN3(n1497), .OUT(n1513) );
  NAND3X1 U1672 ( .IN1(n1502), .IN2(n1501), .IN3(n1500), .OUT(n1504) );
  NOR2X1 U1673 ( .IN1(n1504), .IN2(n1503), .OUT(n1507) );
  NAND3X1 U1674 ( .IN1(n1507), .IN2(n1506), .IN3(n1505), .OUT(n1508) );
  OAI21 U1675 ( .IN1(n1511), .IN2(n1510), .IN3(n414), .OUT(n1512) );
  AOI22 U1676 ( .IN1(Debug_reg[1]), .IN2(n1535), .IN3(n1534), .IN4(n1514), 
        .OUT(n1515) );
  AOI22 U1677 ( .IN1(n1588), .IN2(Debug_reg[1]), .IN3(StateMC[1]), .IN4(n1587), 
        .OUT(n1516) );
  AOI21 U1678 ( .IN1(n1519), .IN2(n1518), .IN3(n1517), .OUT(n1526) );
  NAND3X1 U1679 ( .IN1(n1521), .IN2(n1520), .IN3(n1531), .OUT(n1525) );
  NAND3X1 U1680 ( .IN1(n1526), .IN2(n1525), .IN3(n1524), .OUT(n1527) );
  AOI22 U1681 ( .IN1(Debug_reg[2]), .IN2(n1535), .IN3(n1534), .IN4(n1527), 
        .OUT(n1528) );
  AOI22 U1682 ( .IN1(n1588), .IN2(Debug_reg[2]), .IN3(StateMC[2]), .IN4(n1587), 
        .OUT(n1529) );
  OAI21 U1683 ( .IN1(n1532), .IN2(n1531), .IN3(n1530), .OUT(n1533) );
  AOI22 U1684 ( .IN1(Debug_reg[3]), .IN2(n1535), .IN3(n1534), .IN4(n1533), 
        .OUT(n1536) );
  NOR2X1 U1685 ( .IN1(n317), .IN2(n1539), .OUT(Exc[0]) );
  NOR2X1 U1686 ( .IN1(n223), .IN2(n1539), .OUT(Exc[1]) );
  NOR2X1 U1687 ( .IN1(n222), .IN2(n1539), .OUT(Exc[2]) );
  NOR2X1 U1688 ( .IN1(n308), .IN2(Dataout_valid_BAR), .OUT(Dataout[0]) );
  NOR2X1 U1689 ( .IN1(n298), .IN2(Dataout_valid_BAR), .OUT(Dataout[1]) );
  NOR2X1 U1690 ( .IN1(n311), .IN2(Dataout_valid_BAR), .OUT(Dataout[2]) );
  NOR2X1 U1691 ( .IN1(n186), .IN2(Dataout_valid_BAR), .OUT(Dataout[3]) );
  NOR2X1 U1692 ( .IN1(n309), .IN2(Dataout_valid_BAR), .OUT(Dataout[4]) );
  NOR2X1 U1693 ( .IN1(n314), .IN2(Dataout_valid_BAR), .OUT(Dataout[5]) );
  NOR2X1 U1694 ( .IN1(n310), .IN2(Dataout_valid_BAR), .OUT(Dataout[6]) );
  NOR2X1 U1695 ( .IN1(n396), .IN2(Dataout_valid_BAR), .OUT(Dataout[7]) );
  NOR2X1 U1696 ( .IN1(n406), .IN2(Dataout_valid_BAR), .OUT(Dataout[8]) );
  NOR2X1 U1697 ( .IN1(n293), .IN2(Dataout_valid_BAR), .OUT(Dataout[9]) );
  NOR2X1 U1698 ( .IN1(n294), .IN2(Dataout_valid_BAR), .OUT(Dataout[10]) );
  NOR2X1 U1699 ( .IN1(n408), .IN2(Dataout_valid_BAR), .OUT(Dataout[11]) );
  NOR2X1 U1700 ( .IN1(n304), .IN2(Dataout_valid_BAR), .OUT(Dataout[12]) );
  NOR2X1 U1701 ( .IN1(n295), .IN2(Dataout_valid_BAR), .OUT(Dataout[13]) );
  NOR2X1 U1702 ( .IN1(n405), .IN2(Dataout_valid_BAR), .OUT(Dataout[14]) );
  NOR2X1 U1703 ( .IN1(n1540), .IN2(n1551), .OUT(n1547) );
  OAI21 U1704 ( .IN1(n318), .IN2(n1561), .IN3(n1556), .OUT(n1541) );
  MUX2X1 U1705 ( .IN1(n319), .IN2(add_x_35_A_9_), .S(n1541), .OUT(n1542) );
  NOR2X1 U1706 ( .IN1(n1625), .IN2(n1542), .OUT(n122) );
  MUX2X1 U1707 ( .IN1(n318), .IN2(add_x_35_A_8_), .S(n1543), .OUT(n1544) );
  NOR2X1 U1708 ( .IN1(n1625), .IN2(n1544), .OUT(n121) );
  AOI21 U1709 ( .IN1(n1547), .IN2(add_x_35_A_6_), .IN3(n1548), .OUT(n1545) );
  MUX2X1 U1710 ( .IN1(add_x_35_A_7_), .IN2(n316), .S(n1545), .OUT(n1546) );
  NOR2X1 U1711 ( .IN1(n1625), .IN2(n1546), .OUT(n120) );
  NOR2X1 U1712 ( .IN1(n1548), .IN2(n1547), .OUT(n1549) );
  MUX2X1 U1713 ( .IN1(add_x_35_A_6_), .IN2(n315), .S(n1549), .OUT(n1550) );
  NOR2X1 U1714 ( .IN1(n1625), .IN2(n1550), .OUT(n119) );
  OAI21 U1715 ( .IN1(n1552), .IN2(n1551), .IN3(n1556), .OUT(n1553) );
  MUX2X1 U1716 ( .IN1(n1554), .IN2(add_x_35_A_5_), .S(n1553), .OUT(n1555) );
  NOR2X1 U1717 ( .IN1(n1555), .IN2(n1625), .OUT(n118) );
  OAI21 U1718 ( .IN1(n1560), .IN2(n1561), .IN3(n1556), .OUT(n1559) );
  OAI21 U1719 ( .IN1(n321), .IN2(n1559), .IN3(n1557), .OUT(n1558) );
  AOI21 U1720 ( .IN1(n321), .IN2(n1559), .IN3(n1558), .OUT(n123) );
  INVX1 U1721 ( .IN(Exc_value[1]), .OUT(n1573) );
  INVX1 U1722 ( .IN(Exc_value[2]), .OUT(n1571) );
  AOI22 U1723 ( .IN1(Exc_value[2]), .IN2(Exc_value[0]), .IN3(n1573), .IN4(
        n1571), .OUT(n1572) );
  AOI21 U1724 ( .IN1(Exc_value[0]), .IN2(n1573), .IN3(n1572), .OUT(n1575) );
  NOR2X1 U1725 ( .IN1(n1563), .IN2(n1568), .OUT(n1574) );
  OAI21 U1726 ( .IN1(n1577), .IN2(n1575), .IN3(n1574), .OUT(n1576) );
  OAI21 U1727 ( .IN1(n1566), .IN2(n1576), .IN3(n429), .OUT(n915) );
  NOR2X1 U1728 ( .IN1(n415), .IN2(n1569), .OUT(n1578) );
  AOI22 U1729 ( .IN1(StateMC[0]), .IN2(n1579), .IN3(n1565), .IN4(Exc_Ack), 
        .OUT(n1582) );
  NOR2X1 U1730 ( .IN1(StateMC[0]), .IN2(n1580), .OUT(n1591) );
  NAND3X1 U1731 ( .IN1(n1582), .IN2(n1605), .IN3(n1581), .OUT(n1583) );
  OAI21 U1732 ( .IN1(n1584), .IN2(n1583), .IN3(n429), .OUT(n991) );
  NOR2X1 U1733 ( .IN1(n274), .IN2(Dataout_valid_BAR), .OUT(Dataout[15]) );
  INVX1 U1734 ( .IN(Mode[1]), .OUT(n1586) );
  NAND2X1 U1735 ( .IN1(Mode[0]), .IN2(n1586), .OUT(n1585) );
  NOR2X1 U1736 ( .IN1(Mode[2]), .IN2(n1585), .OUT(n1587) );
  NOR2X1 U1737 ( .IN1(Mode[2]), .IN2(n1586), .OUT(n1588) );
  AOI21 U1738 ( .IN1(n1588), .IN2(Debug_valid_reg), .IN3(n1587), .OUT(n1589)
         );
  NOR2X1 U1739 ( .IN1(n217), .IN2(n1625), .OUT(N254) );
  NOR2X1 U1740 ( .IN1(n216), .IN2(n1625), .OUT(N255) );
  NOR2X1 U1741 ( .IN1(n215), .IN2(n1625), .OUT(N256) );
  NOR2X1 U1742 ( .IN1(n214), .IN2(n1625), .OUT(N257) );
  NOR2X1 U1743 ( .IN1(n213), .IN2(n1625), .OUT(N258) );
  NOR2X1 U1744 ( .IN1(n212), .IN2(n1625), .OUT(N259) );
  INVX1 U1745 ( .IN(Data_valid), .OUT(n1590) );
  NAND2X1 U1746 ( .IN1(n1591), .IN2(n1590), .OUT(n1592) );
  AOI21 U1747 ( .IN1(DP_OP_982J1_125_6202_n182), .IN2(n1615), .IN3(
        DP_OP_982J1_125_6202_n181), .OUT(n1604) );
  AOI22 U1748 ( .IN1(DP_OP_982J1_125_6202_n180), .IN2(
        DP_OP_982J1_125_6202_n136), .IN3(DP_OP_982J1_125_6202_n181), .IN4(
        DP_OP_982J1_125_6202_n135), .OUT(n1603) );
  AOI22 U1749 ( .IN1(Datain1[11]), .IN2(DP_OP_981J1_124_6202_n137), .IN3(
        Datain1[12]), .IN4(n206), .OUT(n1601) );
  AOI22 U1750 ( .IN1(Datain2[7]), .IN2(n200), .IN3(Datain2[8]), .IN4(n272), 
        .OUT(n1593) );
  AOI21 U1751 ( .IN1(Datain1[8]), .IN2(DP_OP_981J1_124_6202_n140), .IN3(n1593), 
        .OUT(n1595) );
  NOR2X1 U1752 ( .IN1(n1595), .IN2(DP_OP_982J1_125_6202_n177), .OUT(n1597) );
  NOR2X1 U1753 ( .IN1(Datain1[10]), .IN2(n1570), .OUT(n1594) );
  AOI21 U1754 ( .IN1(DP_OP_982J1_125_6202_n177), .IN2(n1595), .IN3(n1594), 
        .OUT(n1596) );
  OAI21 U1755 ( .IN1(Datain1[9]), .IN2(n1597), .IN3(n1596), .OUT(n1598) );
  OAI21 U1756 ( .IN1(Datain2[10]), .IN2(n259), .IN3(n1598), .OUT(n1599) );
  OAI21 U1757 ( .IN1(Datain1[11]), .IN2(DP_OP_981J1_124_6202_n137), .IN3(n1599), .OUT(n1600) );
  AOI22 U1758 ( .IN1(DP_OP_982J1_125_6202_n182), .IN2(n1615), .IN3(n1601), 
        .IN4(n1600), .OUT(n1602) );
  OAI21 U1759 ( .IN1(n301), .IN2(n1606), .IN3(n429), .OUT(n1607) );
  OAI21 U1760 ( .IN1(n1607), .IN2(n322), .IN3(n1625), .OUT(n1091) );
  AOI22 U1761 ( .IN1(n1564), .IN2(Datain2[0]), .IN3(n197), .IN4(Datain1[0]), 
        .OUT(n1608) );
  AOI22 U1762 ( .IN1(n1564), .IN2(Datain2[1]), .IN3(n197), .IN4(Datain1[1]), 
        .OUT(n1609) );
  AOI22 U1763 ( .IN1(n1564), .IN2(Datain2[2]), .IN3(n197), .IN4(Datain1[2]), 
        .OUT(n1610) );
  OAI21 U1764 ( .IN1(n413), .IN2(n217), .IN3(n1610), .OUT(n1087) );
  AOI22 U1765 ( .IN1(n1564), .IN2(Datain2[3]), .IN3(n197), .IN4(Datain1[3]), 
        .OUT(n1611) );
  OAI21 U1766 ( .IN1(n413), .IN2(n216), .IN3(n1611), .OUT(n1086) );
  AOI22 U1767 ( .IN1(n1564), .IN2(Datain2[4]), .IN3(n197), .IN4(n416), .OUT(
        n1612) );
  OAI21 U1768 ( .IN1(n413), .IN2(n215), .IN3(n1612), .OUT(n1085) );
  AOI22 U1769 ( .IN1(n1564), .IN2(Datain2[5]), .IN3(n197), .IN4(n417), .OUT(
        n1613) );
  OAI21 U1770 ( .IN1(n413), .IN2(n214), .IN3(n1613), .OUT(n1084) );
  AOI22 U1771 ( .IN1(n1564), .IN2(Datain2[6]), .IN3(n197), .IN4(n418), .OUT(
        n1614) );
  OAI21 U1772 ( .IN1(n413), .IN2(n213), .IN3(n1614), .OUT(n1083) );
  AOI21 U1773 ( .IN1(n197), .IN2(n1621), .IN3(n1564), .OUT(n1616) );
  OAI21 U1774 ( .IN1(n413), .IN2(n212), .IN3(n1616), .OUT(n1082) );
  NOR2X1 U1775 ( .IN1(DP_OP_982J1_125_6202_n181), .IN2(
        DP_OP_982J1_125_6202_n182), .OUT(n1617) );
  NAND3X1 U1776 ( .IN1(n1617), .IN2(DP_OP_981J1_124_6202_n137), .IN3(
        DP_OP_981J1_124_6202_n140), .OUT(n1618) );
  NOR2X1 U1777 ( .IN1(Datain2[7]), .IN2(n1618), .OUT(n1620) );
  NOR2X1 U1778 ( .IN1(DP_OP_982J1_125_6202_n177), .IN2(
        DP_OP_982J1_125_6202_n180), .OUT(n1619) );
  OAI21 U1779 ( .IN1(n1627), .IN2(n1624), .IN3(n1623), .OUT(n1060) );
  OAI21 U1780 ( .IN1(n1628), .IN2(n323), .IN3(n1627), .OUT(n103) );
endmodule


module Mul_cntrl ( CLK, Datain1, Datain2, Data_valid, Dataout, Dataout_valid, 
        Exc, Mode, Debug, Multi_datain1, Multi_datain2, Multi_valid, 
        Multi_dataout, Multi_ack, ExcCheck_valid, ExcCheck_Datain, Exc_value, 
        Exc_Ack, RSTn_BAR );
  input [15:0] Datain1;
  input [15:0] Datain2;
  output [15:0] Dataout;
  output [2:0] Exc;
  input [2:0] Mode;
  output [4:0] Debug;
  output [7:0] Multi_datain1;
  output [7:0] Multi_datain2;
  input [15:0] Multi_dataout;
  output [15:0] ExcCheck_Datain;
  input [2:0] Exc_value;
  input CLK, Data_valid, Multi_ack, Exc_Ack, RSTn_BAR;
  output Dataout_valid, Multi_valid, ExcCheck_valid;
  wire   n1081, StateMC_0_, G_reg, T_reg, N70, N72, N360, N365, N366, N367,
         N368, n59, n89, n96, n97, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n179, n180, n203, n205, n206, n215, n216, n363, n405,
         n417, n521, n548, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         C1_DATA1_8, C1_DATA1_5, C1_DATA1_3, C1_DATA1_2, C1_DATA1_1,
         C1_DATA2_8, C1_DATA2_7, C1_DATA2_6, C1_DATA2_4, C1_DATA2_3,
         C1_DATA2_2, C1_DATA2_1, C1_DATA3_7, C1_DATA3_6, C1_DATA3_5,
         C1_DATA3_2, C1_DATA3_1, C1_DATA4_8, C1_DATA4_7, C1_DATA4_6,
         C1_DATA4_5, C1_DATA4_4, C1_DATA4_3, C1_DATA5_8, C1_DATA5_7,
         C1_DATA5_6, C1_DATA5_5, C1_DATA5_4, C1_DATA5_3, C1_DATA5_2,
         C1_DATA5_1, C1_DATA6_8, C1_DATA6_7, C1_DATA6_6, C1_DATA6_5,
         C1_DATA6_4, C1_DATA6_2, C1_DATA7_8, C1_DATA7_7, C1_DATA7_6,
         C1_DATA7_5, C1_DATA7_4, C1_DATA7_3, C1_DATA7_2, C1_DATA8_8,
         C1_DATA8_7, C1_DATA8_6, C1_DATA8_4, C1_DATA8_0, C1_DATA9_8,
         C1_DATA9_7, C1_DATA9_6, C1_DATA9_5, C1_DATA9_4, C1_DATA9_3,
         C1_DATA9_2, C1_DATA9_0, C1_DATA10_8, C1_DATA10_7, C1_DATA10_6,
         C1_DATA10_5, C1_DATA10_4, C1_DATA10_2, C1_DATA11_8, C1_DATA11_7,
         C1_DATA11_6, C1_DATA11_5, C1_DATA11_3, C1_DATA11_2, C1_DATA11_1,
         C1_DATA12_8, C1_DATA12_7, C1_DATA12_6, C1_DATA12_4, C1_DATA12_3,
         C1_DATA13_8, C1_DATA13_7, C1_DATA13_6, C1_DATA13_5, C1_DATA13_4,
         C1_DATA13_3, C1_DATA13_2, C1_DATA13_1, RSOP_340_C1_Z_0,
         DP_OP_269_159_6943_n103, DP_OP_269_159_6943_n102,
         DP_OP_269_159_6943_n101, DP_OP_269_159_6943_n100,
         DP_OP_269_159_6943_n99, DP_OP_269_159_6943_n98,
         DP_OP_269_159_6943_n97, DP_OP_269_159_6943_n96,
         DP_OP_269_159_6943_n95, DP_OP_269_159_6943_n94,
         DP_OP_269_159_6943_n93, DP_OP_269_159_6943_n92,
         DP_OP_269_159_6943_n91, DP_OP_269_159_6943_n90,
         DP_OP_269_159_6943_n85, DP_OP_269_159_6943_n83,
         DP_OP_269_159_6943_n82, DP_OP_269_159_6943_n79,
         DP_OP_269_159_6943_n78, DP_OP_269_159_6943_n77,
         DP_OP_269_159_6943_n76, DP_OP_269_159_6943_n75,
         DP_OP_269_159_6943_n74, DP_OP_269_159_6943_n73,
         DP_OP_269_159_6943_n72, DP_OP_269_159_6943_n71,
         DP_OP_269_159_6943_n70, DP_OP_269_159_6943_n69,
         DP_OP_269_159_6943_n68, DP_OP_269_159_6943_n67,
         DP_OP_269_159_6943_n66, DP_OP_269_159_6943_n65,
         DP_OP_269_159_6943_n64, DP_OP_269_159_6943_n63,
         DP_OP_269_159_6943_n62, DP_OP_269_159_6943_n61,
         DP_OP_269_159_6943_n60, DP_OP_269_159_6943_n58,
         DP_OP_269_159_6943_n57, DP_OP_269_159_6943_n56,
         DP_OP_269_159_6943_n55, DP_OP_269_159_6943_n51,
         DP_OP_269_159_6943_n50, DP_OP_269_159_6943_n49,
         DP_OP_269_159_6943_n48, DP_OP_269_159_6943_n46,
         DP_OP_269_159_6943_n44, DP_OP_269_159_6943_n43,
         DP_OP_269_159_6943_n42, DP_OP_269_159_6943_n41,
         DP_OP_269_159_6943_n40, DP_OP_269_159_6943_n39,
         DP_OP_269_159_6943_n38, DP_OP_269_159_6943_n34,
         DP_OP_269_159_6943_n29, DP_OP_269_159_6943_n4, DP_OP_269_159_6943_n3,
         DP_OP_349_170_2358_n58, DP_OP_349_170_2358_n57,
         DP_OP_349_170_2358_n56, DP_OP_349_170_2358_n55,
         DP_OP_349_170_2358_n36, DP_OP_349_170_2358_n35,
         DP_OP_349_170_2358_n34, DP_OP_349_170_2358_n33,
         DP_OP_349_170_2358_n32, DP_OP_349_170_2358_n27,
         DP_OP_349_170_2358_n25, DP_OP_349_170_2358_n24,
         DP_OP_349_170_2358_n23, DP_OP_349_170_2358_n21,
         DP_OP_349_170_2358_n20, DP_OP_349_170_2358_n19,
         DP_OP_349_170_2358_n15, DP_OP_349_170_2358_n13,
         DP_OP_349_170_2358_n12, DP_OP_349_170_2358_n11, DP_OP_349_170_2358_n9,
         DP_OP_349_170_2358_n8, DP_OP_349_170_2358_n7, DP_OP_349_170_2358_n3,
         DP_OP_349_170_2358_n2, DP_OP_349_170_2358_n1, DP_OP_347_168_2358_n38,
         DP_OP_347_168_2358_n37, DP_OP_347_168_2358_n36,
         DP_OP_347_168_2358_n35, DP_OP_347_168_2358_n34,
         DP_OP_347_168_2358_n33, DP_OP_347_168_2358_n31,
         DP_OP_347_168_2358_n23, DP_OP_347_168_2358_n21,
         DP_OP_347_168_2358_n20, DP_OP_347_168_2358_n19,
         DP_OP_347_168_2358_n15, DP_OP_347_168_2358_n13,
         DP_OP_347_168_2358_n12, DP_OP_347_168_2358_n11, DP_OP_347_168_2358_n7,
         DP_OP_351_172_2358_n36, DP_OP_351_172_2358_n35,
         DP_OP_351_172_2358_n34, DP_OP_351_172_2358_n33,
         DP_OP_351_172_2358_n31, DP_OP_351_172_2358_n29,
         DP_OP_351_172_2358_n28, DP_OP_351_172_2358_n27,
         DP_OP_351_172_2358_n25, DP_OP_351_172_2358_n24,
         DP_OP_351_172_2358_n23, DP_OP_351_172_2358_n21,
         DP_OP_351_172_2358_n20, DP_OP_351_172_2358_n19,
         DP_OP_351_172_2358_n17, DP_OP_351_172_2358_n16,
         DP_OP_351_172_2358_n15, DP_OP_351_172_2358_n13,
         DP_OP_351_172_2358_n12, DP_OP_351_172_2358_n11, DP_OP_351_172_2358_n9,
         DP_OP_351_172_2358_n8, DP_OP_351_172_2358_n7, DP_OP_341_162_2358_n38,
         DP_OP_341_162_2358_n37, DP_OP_341_162_2358_n36,
         DP_OP_341_162_2358_n34, DP_OP_341_162_2358_n33,
         DP_OP_341_162_2358_n29, DP_OP_341_162_2358_n28,
         DP_OP_341_162_2358_n27, DP_OP_341_162_2358_n25,
         DP_OP_341_162_2358_n24, DP_OP_341_162_2358_n23,
         DP_OP_341_162_2358_n19, DP_OP_341_162_2358_n17,
         DP_OP_341_162_2358_n16, DP_OP_341_162_2358_n15,
         DP_OP_341_162_2358_n13, DP_OP_341_162_2358_n12,
         DP_OP_341_162_2358_n11, DP_OP_341_162_2358_n7, DP_OP_341_162_2358_n5,
         DP_OP_341_162_2358_n4, DP_OP_341_162_2358_n3, DP_OP_345_166_2358_n36,
         DP_OP_345_166_2358_n35, DP_OP_345_166_2358_n34,
         DP_OP_345_166_2358_n33, DP_OP_345_166_2358_n31,
         DP_OP_345_166_2358_n23, DP_OP_345_166_2358_n21,
         DP_OP_345_166_2358_n20, DP_OP_345_166_2358_n19,
         DP_OP_345_166_2358_n17, DP_OP_345_166_2358_n16,
         DP_OP_345_166_2358_n15, DP_OP_345_166_2358_n13,
         DP_OP_345_166_2358_n12, DP_OP_345_166_2358_n11, DP_OP_345_166_2358_n7,
         DP_OP_339_160_2358_n37, DP_OP_339_160_2358_n36,
         DP_OP_339_160_2358_n35, DP_OP_339_160_2358_n33,
         DP_OP_339_160_2358_n32, DP_OP_339_160_2358_n27,
         DP_OP_339_160_2358_n25, DP_OP_339_160_2358_n24,
         DP_OP_339_160_2358_n23, DP_OP_339_160_2358_n21,
         DP_OP_339_160_2358_n20, DP_OP_339_160_2358_n19,
         DP_OP_339_160_2358_n15, DP_OP_339_160_2358_n13,
         DP_OP_339_160_2358_n12, DP_OP_339_160_2358_n7, DP_OP_343_164_2358_n38,
         DP_OP_343_164_2358_n37, DP_OP_343_164_2358_n36,
         DP_OP_343_164_2358_n32, DP_OP_343_164_2358_n29,
         DP_OP_343_164_2358_n28, DP_OP_343_164_2358_n27,
         DP_OP_343_164_2358_n25, DP_OP_343_164_2358_n24,
         DP_OP_343_164_2358_n23, DP_OP_343_164_2358_n21,
         DP_OP_343_164_2358_n20, DP_OP_343_164_2358_n15,
         DP_OP_343_164_2358_n13, DP_OP_343_164_2358_n12, DP_OP_343_164_2358_n7,
         DP_OP_343_164_2358_n5, DP_OP_343_164_2358_n4, DP_OP_343_164_2358_n3,
         DP_OP_343_164_2358_n2, DP_OP_343_164_2358_n1, DP_OP_344_165_2358_n33,
         DP_OP_344_165_2358_n32, DP_OP_344_165_2358_n31,
         DP_OP_344_165_2358_n30, DP_OP_344_165_2358_n29,
         DP_OP_344_165_2358_n28, DP_OP_344_165_2358_n23,
         DP_OP_344_165_2358_n19, DP_OP_344_165_2358_n17,
         DP_OP_344_165_2358_n16, DP_OP_344_165_2358_n15,
         DP_OP_344_165_2358_n13, DP_OP_344_165_2358_n12, DP_OP_344_165_2358_n7,
         DP_OP_344_165_2358_n5, DP_OP_344_165_2358_n4, DP_OP_340_161_2358_n32,
         DP_OP_340_161_2358_n31, DP_OP_340_161_2358_n30,
         DP_OP_340_161_2358_n29, DP_OP_340_161_2358_n28,
         DP_OP_340_161_2358_n27, DP_OP_340_161_2358_n25,
         DP_OP_340_161_2358_n24, DP_OP_340_161_2358_n23,
         DP_OP_340_161_2358_n21, DP_OP_340_161_2358_n20,
         DP_OP_340_161_2358_n15, DP_OP_340_161_2358_n11, DP_OP_340_161_2358_n9,
         DP_OP_340_161_2358_n8, DP_OP_340_161_2358_n7, DP_OP_340_161_2358_n5,
         DP_OP_340_161_2358_n4, DP_OP_340_161_2358_n3, DP_OP_340_161_2358_n2,
         DP_OP_340_161_2358_n1, DP_OP_348_169_2358_n32, DP_OP_348_169_2358_n31,
         DP_OP_348_169_2358_n30, DP_OP_348_169_2358_n29,
         DP_OP_348_169_2358_n23, DP_OP_348_169_2358_n19,
         DP_OP_348_169_2358_n17, DP_OP_348_169_2358_n16,
         DP_OP_348_169_2358_n15, DP_OP_348_169_2358_n13,
         DP_OP_348_169_2358_n12, DP_OP_348_169_2358_n11, DP_OP_348_169_2358_n7,
         DP_OP_348_169_2358_n5, DP_OP_348_169_2358_n4, DP_OP_350_171_2358_n28,
         DP_OP_350_171_2358_n27, DP_OP_350_171_2358_n26,
         DP_OP_350_171_2358_n25, DP_OP_350_171_2358_n24,
         DP_OP_350_171_2358_n23, DP_OP_350_171_2358_n19,
         DP_OP_350_171_2358_n17, DP_OP_350_171_2358_n16,
         DP_OP_350_171_2358_n15, DP_OP_350_171_2358_n13,
         DP_OP_350_171_2358_n11, DP_OP_350_171_2358_n7, DP_OP_350_171_2358_n3,
         DP_OP_350_171_2358_n2, DP_OP_350_171_2358_n1, DP_OP_342_163_2358_n28,
         DP_OP_342_163_2358_n26, DP_OP_342_163_2358_n25,
         DP_OP_342_163_2358_n24, DP_OP_342_163_2358_n23,
         DP_OP_342_163_2358_n21, DP_OP_342_163_2358_n20,
         DP_OP_342_163_2358_n15, DP_OP_342_163_2358_n13,
         DP_OP_342_163_2358_n12, DP_OP_342_163_2358_n11, DP_OP_342_163_2358_n9,
         DP_OP_342_163_2358_n8, DP_OP_342_163_2358_n7, DP_OP_342_163_2358_n5,
         DP_OP_342_163_2358_n4, DP_OP_342_163_2358_n3, DP_OP_342_163_2358_n2,
         DP_OP_342_163_2358_n1, DP_OP_346_167_2358_n23, DP_OP_346_167_2358_n22,
         DP_OP_346_167_2358_n21, DP_OP_346_167_2358_n19,
         DP_OP_346_167_2358_n17, DP_OP_346_167_2358_n16,
         DP_OP_346_167_2358_n15, DP_OP_346_167_2358_n11, DP_OP_346_167_2358_n7,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n90, n91, n92, n93, n94, n95, n98, n115, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n174, n175, n176, n177, n178, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n204,
         n207, n208, n209, n210, n211, n212, n213, n214, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n401, n402, n403, n404, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080;
  wire   [7:0] Final_Exponent_reg;
  wire   [7:0] Op1_Mantissa_reg;
  wire   [7:0] Op2_Mantissa_reg;
  wire   [6:0] Final_Mantissa_reg;

  DFFRX1 T_reg_reg ( .D(n96), .CLK(CLK), .CLRB(n59), .Q(T_reg), .QB(n201) );
  DFFRX1 exc_reg_reg_2_ ( .D(n521), .CLK(CLK), .CLRB(n59), .Q(n203), .QB(n193)
         );
  DFFRX1 exc_reg_reg_0_ ( .D(n405), .CLK(CLK), .CLRB(n59), .Q(n206), .QB(n200)
         );
  DFFRX1 StateMC_reg_1_ ( .D(n548), .CLK(CLK), .CLRB(n59), .Q(n180), .QB(n191)
         );
  DFFRX1 exc_reg_reg_1_ ( .D(n417), .CLK(CLK), .CLRB(n59), .Q(n205), .QB(n202)
         );
  DFFRX1 StateMC_reg_2_ ( .D(N72), .CLK(CLK), .CLRB(n59), .Q(n186), .QB(n179)
         );
  DFFRX1 StateMC_reg_0_ ( .D(N70), .CLK(CLK), .CLRB(n59), .Q(StateMC_0_), .QB(
        n192) );
  DFFRX1 Op1_Mantissa_reg_reg_0_ ( .D(n116), .CLK(CLK), .CLRB(n59), .Q(
        Op1_Mantissa_reg[0]) );
  DFFRX1 Op1_Mantissa_reg_reg_1_ ( .D(n117), .CLK(CLK), .CLRB(n59), .Q(
        Op1_Mantissa_reg[1]) );
  DFFRX1 Op1_Mantissa_reg_reg_2_ ( .D(n118), .CLK(CLK), .CLRB(n59), .Q(
        Op1_Mantissa_reg[2]) );
  DFFRX1 Op1_Mantissa_reg_reg_3_ ( .D(n119), .CLK(CLK), .CLRB(n59), .Q(
        Op1_Mantissa_reg[3]) );
  DFFRX1 Op1_Mantissa_reg_reg_4_ ( .D(n120), .CLK(CLK), .CLRB(n59), .Q(
        Op1_Mantissa_reg[4]) );
  DFFRX1 Op1_Mantissa_reg_reg_5_ ( .D(n121), .CLK(CLK), .CLRB(n59), .Q(
        Op1_Mantissa_reg[5]) );
  DFFRX1 Op1_Mantissa_reg_reg_6_ ( .D(n122), .CLK(CLK), .CLRB(n59), .Q(
        Op1_Mantissa_reg[6]) );
  DFFRX1 Op1_Mantissa_reg_reg_7_ ( .D(n123), .CLK(CLK), .CLRB(n59), .Q(
        Op1_Mantissa_reg[7]) );
  DFFRX1 Op2_Mantissa_reg_reg_6_ ( .D(n130), .CLK(CLK), .CLRB(n59), .Q(
        Op2_Mantissa_reg[6]) );
  DFFRX1 Op2_Mantissa_reg_reg_7_ ( .D(n685), .CLK(CLK), .CLRB(n59), .Q(
        Op2_Mantissa_reg[7]), .QB(n204) );
  DFFRX1 Op2_Mantissa_reg_reg_5_ ( .D(n129), .CLK(CLK), .CLRB(n59), .Q(
        Op2_Mantissa_reg[5]) );
  DFFRX1 Op2_Mantissa_reg_reg_4_ ( .D(n128), .CLK(CLK), .CLRB(n59), .Q(
        Op2_Mantissa_reg[4]) );
  DFFRX1 Op2_Mantissa_reg_reg_3_ ( .D(n127), .CLK(CLK), .CLRB(n59), .Q(
        Op2_Mantissa_reg[3]) );
  DFFRX1 Op2_Mantissa_reg_reg_2_ ( .D(n126), .CLK(CLK), .CLRB(n59), .Q(
        Op2_Mantissa_reg[2]) );
  DFFRX1 Op2_Mantissa_reg_reg_1_ ( .D(n125), .CLK(CLK), .CLRB(n59), .Q(
        Op2_Mantissa_reg[1]) );
  DFFRX1 Op2_Mantissa_reg_reg_0_ ( .D(n124), .CLK(CLK), .CLRB(n59), .Q(
        Op2_Mantissa_reg[0]) );
  DFFRX1 Final_Exponent_reg_reg_8_ ( .D(n89), .CLK(CLK), .CLRB(n59), .QB(n189)
         );
  DFFRX1 ExcCheck_valid_reg ( .D(n684), .CLK(CLK), .CLRB(n59), .Q(
        ExcCheck_valid) );
  DFFRX1 Final_Exponent_reg_reg_0_ ( .D(n691), .CLK(CLK), .CLRB(n59), .Q(
        Final_Exponent_reg[0]), .QB(n393) );
  DFFRX1 Final_Exponent_reg_reg_1_ ( .D(n692), .CLK(CLK), .CLRB(n59), .Q(
        Final_Exponent_reg[1]), .QB(n190) );
  DFFRX1 Final_Exponent_reg_reg_2_ ( .D(n693), .CLK(CLK), .CLRB(n59), .Q(
        Final_Exponent_reg[2]), .QB(n166) );
  DFFRX1 Final_Exponent_reg_reg_3_ ( .D(n694), .CLK(CLK), .CLRB(n59), .Q(
        Final_Exponent_reg[3]), .QB(n165) );
  DFFRX1 Final_Mantissa_reg_reg_0_ ( .D(n363), .CLK(CLK), .CLRB(n59), .Q(n196), 
        .QB(Final_Mantissa_reg[0]) );
  DFFRX1 Final_Mantissa_reg_reg_3_ ( .D(n688), .CLK(CLK), .CLRB(n59), .Q(
        Final_Mantissa_reg[3]), .QB(n195) );
  DFFRX1 Final_Mantissa_reg_reg_4_ ( .D(n689), .CLK(CLK), .CLRB(n59), .Q(
        Final_Mantissa_reg[4]), .QB(n187) );
  DFFRX1 Final_Mantissa_reg_reg_5_ ( .D(n690), .CLK(CLK), .CLRB(n59), .Q(
        Final_Mantissa_reg[5]), .QB(n197) );
  DFFRX1 Final_Mantissa_reg_reg_6_ ( .D(n699), .CLK(CLK), .CLRB(n59), .Q(
        Final_Mantissa_reg[6]), .QB(n198) );
  DFFRX1 Final_Mantissa_reg_reg_1_ ( .D(n686), .CLK(CLK), .CLRB(n59), .Q(
        Final_Mantissa_reg[1]), .QB(n199) );
  DFFRX1 Final_Mantissa_reg_reg_2_ ( .D(n687), .CLK(CLK), .CLRB(n59), .Q(
        Final_Mantissa_reg[2]), .QB(n194) );
  DFFRX1 Final_Exponent_reg_reg_4_ ( .D(n695), .CLK(CLK), .CLRB(n59), .Q(
        Final_Exponent_reg[4]), .QB(n183) );
  DFFRX1 Final_Exponent_reg_reg_5_ ( .D(n696), .CLK(CLK), .CLRB(n59), .Q(
        Final_Exponent_reg[5]), .QB(n185) );
  DFFRX1 Final_Exponent_reg_reg_6_ ( .D(n697), .CLK(CLK), .CLRB(n59), .Q(
        Final_Exponent_reg[6]), .QB(n184) );
  DFFRX1 Final_Exponent_reg_reg_7_ ( .D(n698), .CLK(CLK), .CLRB(n59), .Q(
        Final_Exponent_reg[7]), .QB(n178) );
  DFFRX1 G_reg_reg ( .D(n97), .CLK(CLK), .CLRB(n59), .Q(G_reg), .QB(n188) );
  DFFRX1 Final_Sign_reg_reg ( .D(n683), .CLK(CLK), .CLRB(n59), .Q(n207), .QB(
        n215) );
  DFFRX1 Multi_datain1_reg_7_ ( .D(n106), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain1[7]) );
  DFFRX1 Multi_datain1_reg_6_ ( .D(n105), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain1[6]) );
  DFFRX1 Multi_datain1_reg_5_ ( .D(n104), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain1[5]) );
  DFFRX1 Multi_datain1_reg_4_ ( .D(n103), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain1[4]) );
  DFFRX1 Multi_datain1_reg_3_ ( .D(n102), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain1[3]) );
  DFFRX1 Multi_datain1_reg_2_ ( .D(n101), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain1[2]) );
  DFFRX1 Multi_datain1_reg_1_ ( .D(n100), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain1[1]) );
  DFFRX1 Multi_datain1_reg_0_ ( .D(n99), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain1[0]) );
  DFFRX1 Multi_datain2_reg_7_ ( .D(n114), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain2[7]) );
  DFFRX1 Multi_datain2_reg_6_ ( .D(n113), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain2[6]) );
  DFFRX1 Multi_datain2_reg_5_ ( .D(n112), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain2[5]) );
  DFFRX1 Multi_datain2_reg_4_ ( .D(n111), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain2[4]) );
  DFFRX1 Multi_datain2_reg_3_ ( .D(n110), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain2[3]) );
  DFFRX1 Multi_datain2_reg_2_ ( .D(n109), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain2[2]) );
  DFFRX1 Multi_datain2_reg_1_ ( .D(n108), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain2[1]) );
  DFFRX1 Multi_datain2_reg_0_ ( .D(n107), .CLK(CLK), .CLRB(n59), .Q(
        Multi_datain2[0]) );
  DFFRX1 Multi_valid_reg ( .D(n682), .CLK(CLK), .CLRB(n59), .Q(Multi_valid), 
        .QB(n216) );
  NOR2X1 DP_OP_269_159_6943_U100 ( .IN1(Datain1[14]), .IN2(Datain2[14]), .OUT(
        DP_OP_269_159_6943_n90) );
  NAND2X1 DP_OP_269_159_6943_U95 ( .IN1(Datain2[7]), .IN2(Datain1[7]), .OUT(
        DP_OP_269_159_6943_n78) );
  NOR2X1 DP_OP_269_159_6943_U94 ( .IN1(Datain1[7]), .IN2(Datain2[7]), .OUT(
        DP_OP_269_159_6943_n77) );
  AOI21 DP_OP_269_159_6943_U89 ( .IN1(DP_OP_269_159_6943_n75), .IN2(
        RSOP_340_C1_Z_0), .IN3(DP_OP_269_159_6943_n76), .OUT(
        DP_OP_269_159_6943_n74) );
  NOR2X1 DP_OP_269_159_6943_U83 ( .IN1(n431), .IN2(DP_OP_269_159_6943_n103), 
        .OUT(DP_OP_269_159_6943_n72) );
  OAI21 DP_OP_269_159_6943_U80 ( .IN1(DP_OP_269_159_6943_n74), .IN2(
        DP_OP_269_159_6943_n72), .IN3(DP_OP_269_159_6943_n73), .OUT(
        DP_OP_269_159_6943_n71) );
  NOR2X1 DP_OP_269_159_6943_U73 ( .IN1(DP_OP_269_159_6943_n102), .IN2(
        DP_OP_269_159_6943_n101), .OUT(DP_OP_269_159_6943_n68) );
  OAI21 DP_OP_269_159_6943_U70 ( .IN1(DP_OP_269_159_6943_n68), .IN2(
        DP_OP_269_159_6943_n70), .IN3(DP_OP_269_159_6943_n69), .OUT(
        DP_OP_269_159_6943_n67) );
  NOR2X1 DP_OP_269_159_6943_U64 ( .IN1(DP_OP_269_159_6943_n100), .IN2(
        DP_OP_269_159_6943_n99), .OUT(DP_OP_269_159_6943_n65) );
  OAI21 DP_OP_269_159_6943_U61 ( .IN1(DP_OP_269_159_6943_n69), .IN2(
        DP_OP_269_159_6943_n65), .IN3(DP_OP_269_159_6943_n66), .OUT(
        DP_OP_269_159_6943_n64) );
  NOR2X1 DP_OP_269_159_6943_U60 ( .IN1(DP_OP_269_159_6943_n65), .IN2(
        DP_OP_269_159_6943_n68), .OUT(DP_OP_269_159_6943_n63) );
  AOI21 DP_OP_269_159_6943_U59 ( .IN1(DP_OP_269_159_6943_n63), .IN2(
        DP_OP_269_159_6943_n71), .IN3(DP_OP_269_159_6943_n64), .OUT(
        DP_OP_269_159_6943_n62) );
  NOR2X1 DP_OP_269_159_6943_U53 ( .IN1(DP_OP_269_159_6943_n98), .IN2(
        DP_OP_269_159_6943_n97), .OUT(DP_OP_269_159_6943_n60) );
  NOR2X1 DP_OP_269_159_6943_U44 ( .IN1(DP_OP_269_159_6943_n96), .IN2(
        DP_OP_269_159_6943_n95), .OUT(DP_OP_269_159_6943_n57) );
  OAI21 DP_OP_269_159_6943_U41 ( .IN1(DP_OP_269_159_6943_n61), .IN2(
        DP_OP_269_159_6943_n57), .IN3(DP_OP_269_159_6943_n58), .OUT(
        DP_OP_269_159_6943_n56) );
  NOR2X1 DP_OP_269_159_6943_U40 ( .IN1(DP_OP_269_159_6943_n57), .IN2(
        DP_OP_269_159_6943_n60), .OUT(DP_OP_269_159_6943_n55) );
  NOR2X1 DP_OP_269_159_6943_U31 ( .IN1(DP_OP_269_159_6943_n94), .IN2(
        DP_OP_269_159_6943_n93), .OUT(DP_OP_269_159_6943_n50) );
  NAND2X1 DP_OP_269_159_6943_U25 ( .IN1(DP_OP_269_159_6943_n55), .IN2(
        DP_OP_269_159_6943_n48), .OUT(DP_OP_269_159_6943_n46) );
  NOR2X1 DP_OP_269_159_6943_U18 ( .IN1(DP_OP_269_159_6943_n91), .IN2(
        DP_OP_269_159_6943_n92), .OUT(DP_OP_269_159_6943_n43) );
  OAI21 DP_OP_269_159_6943_U15 ( .IN1(DP_OP_269_159_6943_n51), .IN2(
        DP_OP_269_159_6943_n43), .IN3(DP_OP_269_159_6943_n44), .OUT(
        DP_OP_269_159_6943_n42) );
  NOR2X1 DP_OP_269_159_6943_U14 ( .IN1(DP_OP_269_159_6943_n43), .IN2(
        DP_OP_269_159_6943_n50), .OUT(DP_OP_269_159_6943_n41) );
  AOI21 DP_OP_269_159_6943_U13 ( .IN1(DP_OP_269_159_6943_n41), .IN2(
        DP_OP_269_159_6943_n56), .IN3(DP_OP_269_159_6943_n42), .OUT(
        DP_OP_269_159_6943_n40) );
  OAI21 DP_OP_269_159_6943_U11 ( .IN1(DP_OP_269_159_6943_n39), .IN2(
        DP_OP_269_159_6943_n62), .IN3(DP_OP_269_159_6943_n40), .OUT(
        DP_OP_269_159_6943_n38) );
  NOR2X1 DP_OP_269_159_6943_U5 ( .IN1(DP_OP_269_159_6943_n38), .IN2(
        DP_OP_269_159_6943_n29), .OUT(DP_OP_269_159_6943_n4) );
  NOR2X1 DP_OP_269_159_6943_U4 ( .IN1(DP_OP_269_159_6943_n38), .IN2(
        DP_OP_269_159_6943_n4), .OUT(DP_OP_269_159_6943_n3) );
  NOR2X1 DP_OP_349_170_2358_U40 ( .IN1(n394), .IN2(DP_OP_341_162_2358_n38), 
        .OUT(DP_OP_349_170_2358_n27) );
  NOR2X1 DP_OP_349_170_2358_U37 ( .IN1(DP_OP_341_162_2358_n38), .IN2(
        DP_OP_349_170_2358_n27), .OUT(DP_OP_349_170_2358_n25) );
  NOR2X1 DP_OP_349_170_2358_U36 ( .IN1(n394), .IN2(DP_OP_349_170_2358_n27), 
        .OUT(DP_OP_349_170_2358_n24) );
  NOR2X1 DP_OP_349_170_2358_U35 ( .IN1(DP_OP_349_170_2358_n25), .IN2(
        DP_OP_349_170_2358_n24), .OUT(C1_DATA11_2) );
  NOR2X1 DP_OP_349_170_2358_U19 ( .IN1(DP_OP_349_170_2358_n35), .IN2(
        DP_OP_349_170_2358_n15), .OUT(DP_OP_349_170_2358_n13) );
  NOR2X1 DP_OP_349_170_2358_U18 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_349_170_2358_n15), .OUT(DP_OP_349_170_2358_n12) );
  NOR2X1 DP_OP_349_170_2358_U17 ( .IN1(DP_OP_349_170_2358_n13), .IN2(
        DP_OP_349_170_2358_n12), .OUT(C1_DATA11_5) );
  NOR2X1 DP_OP_349_170_2358_U16 ( .IN1(DP_OP_349_170_2358_n58), .IN2(
        DP_OP_349_170_2358_n34), .OUT(DP_OP_349_170_2358_n11) );
  NOR2X1 DP_OP_349_170_2358_U13 ( .IN1(DP_OP_349_170_2358_n34), .IN2(
        DP_OP_349_170_2358_n11), .OUT(DP_OP_349_170_2358_n9) );
  NOR2X1 DP_OP_349_170_2358_U12 ( .IN1(DP_OP_349_170_2358_n58), .IN2(
        DP_OP_349_170_2358_n11), .OUT(DP_OP_349_170_2358_n8) );
  NOR2X1 DP_OP_349_170_2358_U11 ( .IN1(DP_OP_349_170_2358_n9), .IN2(
        DP_OP_349_170_2358_n8), .OUT(C1_DATA11_6) );
  NOR2X1 DP_OP_349_170_2358_U10 ( .IN1(n181), .IN2(DP_OP_349_170_2358_n33), 
        .OUT(DP_OP_349_170_2358_n7) );
  NOR2X1 DP_OP_349_170_2358_U4 ( .IN1(DP_OP_349_170_2358_n32), .IN2(n408), 
        .OUT(DP_OP_349_170_2358_n3) );
  NOR2X1 DP_OP_349_170_2358_U3 ( .IN1(DP_OP_349_170_2358_n32), .IN2(
        DP_OP_349_170_2358_n3), .OUT(DP_OP_349_170_2358_n2) );
  NOR2X1 DP_OP_349_170_2358_U2 ( .IN1(n408), .IN2(DP_OP_349_170_2358_n3), 
        .OUT(DP_OP_349_170_2358_n1) );
  NOR2X1 DP_OP_349_170_2358_U1 ( .IN1(DP_OP_349_170_2358_n2), .IN2(
        DP_OP_349_170_2358_n1), .OUT(C1_DATA11_8) );
  NOR2X1 DP_OP_347_168_2358_U28 ( .IN1(DP_OP_349_170_2358_n56), .IN2(
        DP_OP_347_168_2358_n36), .OUT(DP_OP_347_168_2358_n19) );
  NOR2X1 DP_OP_347_168_2358_U22 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_347_168_2358_n35), .OUT(DP_OP_347_168_2358_n15) );
  NOR2X1 DP_OP_347_168_2358_U19 ( .IN1(DP_OP_347_168_2358_n35), .IN2(
        DP_OP_347_168_2358_n15), .OUT(DP_OP_347_168_2358_n13) );
  NOR2X1 DP_OP_347_168_2358_U18 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_347_168_2358_n15), .OUT(DP_OP_347_168_2358_n12) );
  NOR2X1 DP_OP_347_168_2358_U17 ( .IN1(DP_OP_347_168_2358_n13), .IN2(
        DP_OP_347_168_2358_n12), .OUT(C1_DATA9_5) );
  NOR2X1 DP_OP_347_168_2358_U16 ( .IN1(DP_OP_349_170_2358_n58), .IN2(
        DP_OP_347_168_2358_n34), .OUT(DP_OP_347_168_2358_n11) );
  NOR2X1 DP_OP_347_168_2358_U10 ( .IN1(n181), .IN2(DP_OP_347_168_2358_n33), 
        .OUT(DP_OP_347_168_2358_n7) );
  NOR2X1 DP_OP_351_172_2358_U46 ( .IN1(Final_Exponent_reg[1]), .IN2(
        Final_Exponent_reg[0]), .OUT(DP_OP_351_172_2358_n31) );
  NOR2X1 DP_OP_351_172_2358_U43 ( .IN1(C1_DATA8_0), .IN2(n169), .OUT(
        DP_OP_351_172_2358_n29) );
  NOR2X1 DP_OP_351_172_2358_U42 ( .IN1(n404), .IN2(n169), .OUT(
        DP_OP_351_172_2358_n28) );
  NOR2X1 DP_OP_351_172_2358_U41 ( .IN1(DP_OP_351_172_2358_n29), .IN2(
        DP_OP_351_172_2358_n28), .OUT(C1_DATA13_1) );
  NOR2X1 DP_OP_351_172_2358_U25 ( .IN1(DP_OP_351_172_2358_n36), .IN2(
        DP_OP_351_172_2358_n19), .OUT(DP_OP_351_172_2358_n17) );
  NOR2X1 DP_OP_351_172_2358_U24 ( .IN1(DP_OP_349_170_2358_n56), .IN2(
        DP_OP_351_172_2358_n19), .OUT(DP_OP_351_172_2358_n16) );
  NOR2X1 DP_OP_351_172_2358_U23 ( .IN1(DP_OP_351_172_2358_n17), .IN2(
        DP_OP_351_172_2358_n16), .OUT(C1_DATA13_4) );
  NOR2X1 DP_OP_351_172_2358_U19 ( .IN1(DP_OP_351_172_2358_n35), .IN2(
        DP_OP_351_172_2358_n15), .OUT(DP_OP_351_172_2358_n13) );
  NOR2X1 DP_OP_351_172_2358_U18 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_351_172_2358_n15), .OUT(DP_OP_351_172_2358_n12) );
  NOR2X1 DP_OP_351_172_2358_U17 ( .IN1(DP_OP_351_172_2358_n13), .IN2(
        DP_OP_351_172_2358_n12), .OUT(C1_DATA13_5) );
  NOR2X1 DP_OP_351_172_2358_U16 ( .IN1(DP_OP_349_170_2358_n58), .IN2(
        DP_OP_351_172_2358_n34), .OUT(DP_OP_351_172_2358_n11) );
  NOR2X1 DP_OP_351_172_2358_U13 ( .IN1(DP_OP_351_172_2358_n34), .IN2(
        DP_OP_351_172_2358_n11), .OUT(DP_OP_351_172_2358_n9) );
  NOR2X1 DP_OP_351_172_2358_U12 ( .IN1(DP_OP_349_170_2358_n58), .IN2(
        DP_OP_351_172_2358_n11), .OUT(DP_OP_351_172_2358_n8) );
  NOR2X1 DP_OP_351_172_2358_U11 ( .IN1(DP_OP_351_172_2358_n9), .IN2(
        DP_OP_351_172_2358_n8), .OUT(C1_DATA13_6) );
  NOR2X1 DP_OP_351_172_2358_U10 ( .IN1(n181), .IN2(DP_OP_351_172_2358_n33), 
        .OUT(DP_OP_351_172_2358_n7) );
  NOR2X1 DP_OP_341_162_2358_U40 ( .IN1(Final_Exponent_reg[2]), .IN2(
        DP_OP_341_162_2358_n38), .OUT(DP_OP_341_162_2358_n27) );
  NOR2X1 DP_OP_341_162_2358_U37 ( .IN1(DP_OP_341_162_2358_n38), .IN2(
        DP_OP_341_162_2358_n27), .OUT(DP_OP_341_162_2358_n25) );
  NOR2X1 DP_OP_341_162_2358_U36 ( .IN1(n394), .IN2(DP_OP_341_162_2358_n27), 
        .OUT(DP_OP_341_162_2358_n24) );
  NOR2X1 DP_OP_341_162_2358_U35 ( .IN1(DP_OP_341_162_2358_n25), .IN2(
        DP_OP_341_162_2358_n24), .OUT(C1_DATA3_2) );
  NOR2X1 DP_OP_341_162_2358_U34 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_341_162_2358_n37), .OUT(DP_OP_341_162_2358_n23) );
  NOR2X1 DP_OP_341_162_2358_U25 ( .IN1(DP_OP_341_162_2358_n36), .IN2(
        DP_OP_341_162_2358_n19), .OUT(DP_OP_341_162_2358_n17) );
  NOR2X1 DP_OP_341_162_2358_U24 ( .IN1(DP_OP_349_170_2358_n56), .IN2(
        DP_OP_341_162_2358_n19), .OUT(DP_OP_341_162_2358_n16) );
  NOR2X1 DP_OP_341_162_2358_U22 ( .IN1(DP_OP_349_170_2358_n57), .IN2(n167), 
        .OUT(DP_OP_341_162_2358_n15) );
  NOR2X1 DP_OP_341_162_2358_U19 ( .IN1(n167), .IN2(DP_OP_341_162_2358_n15), 
        .OUT(DP_OP_341_162_2358_n13) );
  NOR2X1 DP_OP_341_162_2358_U18 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_341_162_2358_n15), .OUT(DP_OP_341_162_2358_n12) );
  NOR2X1 DP_OP_341_162_2358_U17 ( .IN1(DP_OP_341_162_2358_n13), .IN2(
        DP_OP_341_162_2358_n12), .OUT(C1_DATA3_5) );
  NOR2X1 DP_OP_341_162_2358_U16 ( .IN1(DP_OP_349_170_2358_n58), .IN2(
        DP_OP_341_162_2358_n34), .OUT(DP_OP_341_162_2358_n11) );
  NOR2X1 DP_OP_341_162_2358_U7 ( .IN1(DP_OP_341_162_2358_n33), .IN2(
        DP_OP_341_162_2358_n7), .OUT(DP_OP_341_162_2358_n5) );
  NOR2X1 DP_OP_341_162_2358_U6 ( .IN1(n181), .IN2(DP_OP_341_162_2358_n7), 
        .OUT(DP_OP_341_162_2358_n4) );
  NOR2X1 DP_OP_341_162_2358_U5 ( .IN1(DP_OP_341_162_2358_n5), .IN2(
        DP_OP_341_162_2358_n4), .OUT(C1_DATA3_7) );
  NOR2X1 DP_OP_341_162_2358_U4 ( .IN1(n177), .IN2(n408), .OUT(
        DP_OP_341_162_2358_n3) );
  NOR2X1 DP_OP_345_166_2358_U31 ( .IN1(n650), .IN2(DP_OP_345_166_2358_n23), 
        .OUT(DP_OP_345_166_2358_n21) );
  NOR2X1 DP_OP_345_166_2358_U30 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_345_166_2358_n23), .OUT(DP_OP_345_166_2358_n20) );
  NOR2X1 DP_OP_345_166_2358_U29 ( .IN1(DP_OP_345_166_2358_n21), .IN2(
        DP_OP_345_166_2358_n20), .OUT(C1_DATA7_3) );
  NOR2X1 DP_OP_345_166_2358_U25 ( .IN1(DP_OP_345_166_2358_n36), .IN2(
        DP_OP_345_166_2358_n19), .OUT(DP_OP_345_166_2358_n17) );
  NOR2X1 DP_OP_345_166_2358_U24 ( .IN1(DP_OP_349_170_2358_n56), .IN2(
        DP_OP_345_166_2358_n19), .OUT(DP_OP_345_166_2358_n16) );
  NOR2X1 DP_OP_345_166_2358_U23 ( .IN1(DP_OP_345_166_2358_n17), .IN2(
        DP_OP_345_166_2358_n16), .OUT(C1_DATA7_4) );
  NOR2X1 DP_OP_345_166_2358_U22 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_345_166_2358_n35), .OUT(DP_OP_345_166_2358_n15) );
  NOR2X1 DP_OP_345_166_2358_U19 ( .IN1(DP_OP_345_166_2358_n35), .IN2(
        DP_OP_345_166_2358_n15), .OUT(DP_OP_345_166_2358_n13) );
  NOR2X1 DP_OP_345_166_2358_U18 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_345_166_2358_n15), .OUT(DP_OP_345_166_2358_n12) );
  NOR2X1 DP_OP_345_166_2358_U17 ( .IN1(DP_OP_345_166_2358_n13), .IN2(
        DP_OP_345_166_2358_n12), .OUT(C1_DATA7_5) );
  NOR2X1 DP_OP_345_166_2358_U16 ( .IN1(DP_OP_349_170_2358_n58), .IN2(
        DP_OP_345_166_2358_n34), .OUT(DP_OP_345_166_2358_n11) );
  NOR2X1 DP_OP_345_166_2358_U10 ( .IN1(n181), .IN2(DP_OP_345_166_2358_n33), 
        .OUT(DP_OP_345_166_2358_n7) );
  NOR2X1 DP_OP_339_160_2358_U41 ( .IN1(DP_OP_351_172_2358_n29), .IN2(
        DP_OP_351_172_2358_n28), .OUT(C1_DATA1_1) );
  NOR2X1 DP_OP_339_160_2358_U40 ( .IN1(Final_Exponent_reg[2]), .IN2(
        DP_OP_343_164_2358_n38), .OUT(DP_OP_339_160_2358_n27) );
  NOR2X1 DP_OP_339_160_2358_U37 ( .IN1(DP_OP_343_164_2358_n38), .IN2(
        DP_OP_339_160_2358_n27), .OUT(DP_OP_339_160_2358_n25) );
  NOR2X1 DP_OP_339_160_2358_U36 ( .IN1(Final_Exponent_reg[2]), .IN2(
        DP_OP_339_160_2358_n27), .OUT(DP_OP_339_160_2358_n24) );
  NOR2X1 DP_OP_339_160_2358_U35 ( .IN1(DP_OP_339_160_2358_n25), .IN2(
        DP_OP_339_160_2358_n24), .OUT(C1_DATA1_2) );
  NOR2X1 DP_OP_339_160_2358_U34 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_339_160_2358_n37), .OUT(DP_OP_339_160_2358_n23) );
  NOR2X1 DP_OP_339_160_2358_U31 ( .IN1(DP_OP_339_160_2358_n37), .IN2(
        DP_OP_339_160_2358_n23), .OUT(DP_OP_339_160_2358_n21) );
  NOR2X1 DP_OP_339_160_2358_U30 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_339_160_2358_n23), .OUT(DP_OP_339_160_2358_n20) );
  NOR2X1 DP_OP_339_160_2358_U29 ( .IN1(DP_OP_339_160_2358_n21), .IN2(
        DP_OP_339_160_2358_n20), .OUT(C1_DATA1_3) );
  NOR2X1 DP_OP_339_160_2358_U28 ( .IN1(DP_OP_349_170_2358_n56), .IN2(
        DP_OP_339_160_2358_n36), .OUT(DP_OP_339_160_2358_n19) );
  NOR2X1 DP_OP_339_160_2358_U22 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_339_160_2358_n35), .OUT(DP_OP_339_160_2358_n15) );
  NOR2X1 DP_OP_339_160_2358_U19 ( .IN1(DP_OP_339_160_2358_n35), .IN2(
        DP_OP_339_160_2358_n15), .OUT(DP_OP_339_160_2358_n13) );
  NOR2X1 DP_OP_339_160_2358_U18 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_339_160_2358_n15), .OUT(DP_OP_339_160_2358_n12) );
  NOR2X1 DP_OP_339_160_2358_U17 ( .IN1(DP_OP_339_160_2358_n13), .IN2(
        DP_OP_339_160_2358_n12), .OUT(C1_DATA1_5) );
  NOR2X1 DP_OP_343_164_2358_U43 ( .IN1(C1_DATA8_0), .IN2(
        DP_OP_351_172_2358_n31), .OUT(DP_OP_343_164_2358_n29) );
  NOR2X1 DP_OP_343_164_2358_U42 ( .IN1(n404), .IN2(DP_OP_351_172_2358_n31), 
        .OUT(DP_OP_343_164_2358_n28) );
  NOR2X1 DP_OP_343_164_2358_U41 ( .IN1(DP_OP_343_164_2358_n29), .IN2(
        DP_OP_343_164_2358_n28), .OUT(C1_DATA5_1) );
  NOR2X1 DP_OP_343_164_2358_U34 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_343_164_2358_n37), .OUT(DP_OP_343_164_2358_n23) );
  NOR2X1 DP_OP_343_164_2358_U31 ( .IN1(DP_OP_343_164_2358_n37), .IN2(n176), 
        .OUT(DP_OP_343_164_2358_n21) );
  NOR2X1 DP_OP_343_164_2358_U30 ( .IN1(DP_OP_349_170_2358_n55), .IN2(n176), 
        .OUT(DP_OP_343_164_2358_n20) );
  NOR2X1 DP_OP_343_164_2358_U29 ( .IN1(DP_OP_343_164_2358_n21), .IN2(
        DP_OP_343_164_2358_n20), .OUT(C1_DATA5_3) );
  NOR2X1 DP_OP_343_164_2358_U22 ( .IN1(DP_OP_349_170_2358_n57), .IN2(n398), 
        .OUT(DP_OP_343_164_2358_n15) );
  NOR2X1 DP_OP_343_164_2358_U19 ( .IN1(n398), .IN2(DP_OP_343_164_2358_n15), 
        .OUT(DP_OP_343_164_2358_n13) );
  NOR2X1 DP_OP_343_164_2358_U18 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_343_164_2358_n15), .OUT(DP_OP_343_164_2358_n12) );
  NOR2X1 DP_OP_343_164_2358_U17 ( .IN1(DP_OP_343_164_2358_n13), .IN2(
        DP_OP_343_164_2358_n12), .OUT(C1_DATA5_5) );
  NOR2X1 DP_OP_343_164_2358_U10 ( .IN1(n181), .IN2(n162), .OUT(
        DP_OP_343_164_2358_n7) );
  NOR2X1 DP_OP_343_164_2358_U7 ( .IN1(n162), .IN2(DP_OP_343_164_2358_n7), 
        .OUT(DP_OP_343_164_2358_n5) );
  NOR2X1 DP_OP_343_164_2358_U6 ( .IN1(n181), .IN2(DP_OP_343_164_2358_n7), 
        .OUT(DP_OP_343_164_2358_n4) );
  NOR2X1 DP_OP_343_164_2358_U5 ( .IN1(DP_OP_343_164_2358_n5), .IN2(
        DP_OP_343_164_2358_n4), .OUT(C1_DATA5_7) );
  NOR2X1 DP_OP_343_164_2358_U4 ( .IN1(DP_OP_343_164_2358_n32), .IN2(n408), 
        .OUT(DP_OP_343_164_2358_n3) );
  NOR2X1 DP_OP_343_164_2358_U3 ( .IN1(DP_OP_343_164_2358_n32), .IN2(
        DP_OP_343_164_2358_n3), .OUT(DP_OP_343_164_2358_n2) );
  NOR2X1 DP_OP_343_164_2358_U2 ( .IN1(n408), .IN2(DP_OP_343_164_2358_n3), 
        .OUT(DP_OP_343_164_2358_n1) );
  NOR2X1 DP_OP_343_164_2358_U1 ( .IN1(DP_OP_343_164_2358_n2), .IN2(
        DP_OP_343_164_2358_n1), .OUT(C1_DATA5_8) );
  NOR2X1 DP_OP_344_165_2358_U34 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_344_165_2358_n33), .OUT(DP_OP_344_165_2358_n23) );
  NOR2X1 DP_OP_344_165_2358_U28 ( .IN1(DP_OP_349_170_2358_n56), .IN2(
        DP_OP_344_165_2358_n32), .OUT(DP_OP_344_165_2358_n19) );
  NOR2X1 DP_OP_344_165_2358_U25 ( .IN1(DP_OP_344_165_2358_n32), .IN2(
        DP_OP_344_165_2358_n19), .OUT(DP_OP_344_165_2358_n17) );
  NOR2X1 DP_OP_344_165_2358_U24 ( .IN1(DP_OP_349_170_2358_n56), .IN2(
        DP_OP_344_165_2358_n19), .OUT(DP_OP_344_165_2358_n16) );
  NOR2X1 DP_OP_344_165_2358_U23 ( .IN1(DP_OP_344_165_2358_n17), .IN2(
        DP_OP_344_165_2358_n16), .OUT(C1_DATA6_4) );
  NOR2X1 DP_OP_344_165_2358_U19 ( .IN1(DP_OP_344_165_2358_n31), .IN2(
        DP_OP_344_165_2358_n15), .OUT(DP_OP_344_165_2358_n13) );
  NOR2X1 DP_OP_344_165_2358_U18 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_344_165_2358_n15), .OUT(DP_OP_344_165_2358_n12) );
  NOR2X1 DP_OP_344_165_2358_U17 ( .IN1(DP_OP_344_165_2358_n13), .IN2(
        DP_OP_344_165_2358_n12), .OUT(C1_DATA6_5) );
  NOR2X1 DP_OP_344_165_2358_U10 ( .IN1(n181), .IN2(DP_OP_344_165_2358_n29), 
        .OUT(DP_OP_344_165_2358_n7) );
  NOR2X1 DP_OP_344_165_2358_U7 ( .IN1(DP_OP_344_165_2358_n29), .IN2(
        DP_OP_344_165_2358_n7), .OUT(DP_OP_344_165_2358_n5) );
  NOR2X1 DP_OP_344_165_2358_U6 ( .IN1(n181), .IN2(DP_OP_344_165_2358_n7), 
        .OUT(DP_OP_344_165_2358_n4) );
  NOR2X1 DP_OP_344_165_2358_U5 ( .IN1(DP_OP_344_165_2358_n5), .IN2(
        DP_OP_344_165_2358_n4), .OUT(C1_DATA6_7) );
  NOR2X1 DP_OP_340_161_2358_U40 ( .IN1(Final_Exponent_reg[2]), .IN2(
        Final_Exponent_reg[1]), .OUT(DP_OP_340_161_2358_n27) );
  NOR2X1 DP_OP_340_161_2358_U37 ( .IN1(n404), .IN2(DP_OP_340_161_2358_n27), 
        .OUT(DP_OP_340_161_2358_n25) );
  NOR2X1 DP_OP_340_161_2358_U36 ( .IN1(n394), .IN2(DP_OP_340_161_2358_n27), 
        .OUT(DP_OP_340_161_2358_n24) );
  NOR2X1 DP_OP_340_161_2358_U35 ( .IN1(DP_OP_340_161_2358_n25), .IN2(
        DP_OP_340_161_2358_n24), .OUT(C1_DATA2_2) );
  NOR2X1 DP_OP_340_161_2358_U31 ( .IN1(n174), .IN2(DP_OP_340_161_2358_n23), 
        .OUT(DP_OP_340_161_2358_n21) );
  NOR2X1 DP_OP_340_161_2358_U30 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_340_161_2358_n23), .OUT(DP_OP_340_161_2358_n20) );
  NOR2X1 DP_OP_340_161_2358_U29 ( .IN1(DP_OP_340_161_2358_n21), .IN2(
        DP_OP_340_161_2358_n20), .OUT(C1_DATA2_3) );
  NOR2X1 DP_OP_340_161_2358_U22 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_340_161_2358_n31), .OUT(DP_OP_340_161_2358_n15) );
  NOR2X1 DP_OP_340_161_2358_U16 ( .IN1(DP_OP_349_170_2358_n58), .IN2(
        DP_OP_340_161_2358_n30), .OUT(DP_OP_340_161_2358_n11) );
  NOR2X1 DP_OP_340_161_2358_U13 ( .IN1(DP_OP_340_161_2358_n30), .IN2(
        DP_OP_340_161_2358_n11), .OUT(DP_OP_340_161_2358_n9) );
  NOR2X1 DP_OP_340_161_2358_U12 ( .IN1(DP_OP_349_170_2358_n58), .IN2(
        DP_OP_340_161_2358_n11), .OUT(DP_OP_340_161_2358_n8) );
  NOR2X1 DP_OP_340_161_2358_U11 ( .IN1(DP_OP_340_161_2358_n9), .IN2(
        DP_OP_340_161_2358_n8), .OUT(C1_DATA2_6) );
  NOR2X1 DP_OP_340_161_2358_U10 ( .IN1(n181), .IN2(DP_OP_340_161_2358_n29), 
        .OUT(DP_OP_340_161_2358_n7) );
  NOR2X1 DP_OP_340_161_2358_U7 ( .IN1(DP_OP_340_161_2358_n29), .IN2(
        DP_OP_340_161_2358_n7), .OUT(DP_OP_340_161_2358_n5) );
  NOR2X1 DP_OP_340_161_2358_U6 ( .IN1(n181), .IN2(DP_OP_340_161_2358_n7), 
        .OUT(DP_OP_340_161_2358_n4) );
  NOR2X1 DP_OP_340_161_2358_U5 ( .IN1(DP_OP_340_161_2358_n5), .IN2(
        DP_OP_340_161_2358_n4), .OUT(C1_DATA2_7) );
  NOR2X1 DP_OP_340_161_2358_U4 ( .IN1(DP_OP_340_161_2358_n28), .IN2(n408), 
        .OUT(DP_OP_340_161_2358_n3) );
  NOR2X1 DP_OP_340_161_2358_U3 ( .IN1(DP_OP_340_161_2358_n28), .IN2(
        DP_OP_340_161_2358_n3), .OUT(DP_OP_340_161_2358_n2) );
  NOR2X1 DP_OP_340_161_2358_U2 ( .IN1(n408), .IN2(DP_OP_340_161_2358_n3), 
        .OUT(DP_OP_340_161_2358_n1) );
  NOR2X1 DP_OP_340_161_2358_U1 ( .IN1(DP_OP_340_161_2358_n2), .IN2(
        DP_OP_340_161_2358_n1), .OUT(C1_DATA2_8) );
  NOR2X1 DP_OP_348_169_2358_U35 ( .IN1(DP_OP_340_161_2358_n25), .IN2(
        DP_OP_340_161_2358_n24), .OUT(C1_DATA10_2) );
  NOR2X1 DP_OP_348_169_2358_U25 ( .IN1(DP_OP_348_169_2358_n32), .IN2(
        DP_OP_348_169_2358_n19), .OUT(DP_OP_348_169_2358_n17) );
  NOR2X1 DP_OP_348_169_2358_U24 ( .IN1(DP_OP_349_170_2358_n56), .IN2(
        DP_OP_348_169_2358_n19), .OUT(DP_OP_348_169_2358_n16) );
  NOR2X1 DP_OP_348_169_2358_U23 ( .IN1(DP_OP_348_169_2358_n17), .IN2(
        DP_OP_348_169_2358_n16), .OUT(C1_DATA10_4) );
  NOR2X1 DP_OP_348_169_2358_U22 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_348_169_2358_n31), .OUT(DP_OP_348_169_2358_n15) );
  NOR2X1 DP_OP_348_169_2358_U19 ( .IN1(DP_OP_348_169_2358_n31), .IN2(
        DP_OP_348_169_2358_n15), .OUT(DP_OP_348_169_2358_n13) );
  NOR2X1 DP_OP_348_169_2358_U18 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_348_169_2358_n15), .OUT(DP_OP_348_169_2358_n12) );
  NOR2X1 DP_OP_348_169_2358_U17 ( .IN1(DP_OP_348_169_2358_n13), .IN2(
        DP_OP_348_169_2358_n12), .OUT(C1_DATA10_5) );
  NOR2X1 DP_OP_348_169_2358_U16 ( .IN1(DP_OP_349_170_2358_n58), .IN2(
        DP_OP_348_169_2358_n30), .OUT(DP_OP_348_169_2358_n11) );
  NOR2X1 DP_OP_348_169_2358_U10 ( .IN1(n181), .IN2(DP_OP_348_169_2358_n29), 
        .OUT(DP_OP_348_169_2358_n7) );
  NOR2X1 DP_OP_348_169_2358_U7 ( .IN1(DP_OP_348_169_2358_n29), .IN2(
        DP_OP_348_169_2358_n7), .OUT(DP_OP_348_169_2358_n5) );
  NOR2X1 DP_OP_348_169_2358_U6 ( .IN1(n181), .IN2(DP_OP_348_169_2358_n7), 
        .OUT(DP_OP_348_169_2358_n4) );
  NOR2X1 DP_OP_348_169_2358_U5 ( .IN1(DP_OP_348_169_2358_n5), .IN2(
        DP_OP_348_169_2358_n4), .OUT(C1_DATA10_7) );
  NOR2X1 DP_OP_350_171_2358_U28 ( .IN1(DP_OP_349_170_2358_n56), .IN2(
        DP_OP_350_171_2358_n28), .OUT(DP_OP_350_171_2358_n19) );
  NOR2X1 DP_OP_350_171_2358_U25 ( .IN1(DP_OP_350_171_2358_n28), .IN2(
        DP_OP_350_171_2358_n19), .OUT(DP_OP_350_171_2358_n17) );
  NOR2X1 DP_OP_350_171_2358_U24 ( .IN1(DP_OP_349_170_2358_n56), .IN2(
        DP_OP_350_171_2358_n19), .OUT(DP_OP_350_171_2358_n16) );
  NOR2X1 DP_OP_350_171_2358_U23 ( .IN1(DP_OP_350_171_2358_n17), .IN2(
        DP_OP_350_171_2358_n16), .OUT(C1_DATA12_4) );
  NOR2X1 DP_OP_350_171_2358_U22 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_350_171_2358_n27), .OUT(DP_OP_350_171_2358_n15) );
  NOR2X1 DP_OP_350_171_2358_U19 ( .IN1(DP_OP_350_171_2358_n27), .IN2(
        DP_OP_350_171_2358_n15), .OUT(DP_OP_350_171_2358_n13) );
  NOR2X1 DP_OP_350_171_2358_U16 ( .IN1(DP_OP_349_170_2358_n58), .IN2(
        DP_OP_350_171_2358_n26), .OUT(DP_OP_350_171_2358_n11) );
  NOR2X1 DP_OP_350_171_2358_U10 ( .IN1(n181), .IN2(DP_OP_350_171_2358_n25), 
        .OUT(DP_OP_350_171_2358_n7) );
  NOR2X1 DP_OP_350_171_2358_U4 ( .IN1(DP_OP_350_171_2358_n24), .IN2(n408), 
        .OUT(DP_OP_350_171_2358_n3) );
  NOR2X1 DP_OP_350_171_2358_U3 ( .IN1(DP_OP_350_171_2358_n24), .IN2(
        DP_OP_350_171_2358_n3), .OUT(DP_OP_350_171_2358_n2) );
  NOR2X1 DP_OP_350_171_2358_U2 ( .IN1(n408), .IN2(DP_OP_350_171_2358_n3), 
        .OUT(DP_OP_350_171_2358_n1) );
  NOR2X1 DP_OP_350_171_2358_U1 ( .IN1(DP_OP_350_171_2358_n2), .IN2(
        DP_OP_350_171_2358_n1), .OUT(C1_DATA12_8) );
  NOR2X1 DP_OP_342_163_2358_U31 ( .IN1(n394), .IN2(DP_OP_342_163_2358_n23), 
        .OUT(DP_OP_342_163_2358_n21) );
  NOR2X1 DP_OP_342_163_2358_U30 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_342_163_2358_n23), .OUT(DP_OP_342_163_2358_n20) );
  NOR2X1 DP_OP_342_163_2358_U29 ( .IN1(DP_OP_342_163_2358_n21), .IN2(
        DP_OP_342_163_2358_n20), .OUT(C1_DATA4_3) );
  NOR2X1 DP_OP_342_163_2358_U22 ( .IN1(DP_OP_349_170_2358_n57), .IN2(n382), 
        .OUT(DP_OP_342_163_2358_n15) );
  NOR2X1 DP_OP_342_163_2358_U19 ( .IN1(n382), .IN2(DP_OP_342_163_2358_n15), 
        .OUT(DP_OP_342_163_2358_n13) );
  NOR2X1 DP_OP_342_163_2358_U18 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_342_163_2358_n15), .OUT(DP_OP_342_163_2358_n12) );
  NOR2X1 DP_OP_342_163_2358_U17 ( .IN1(DP_OP_342_163_2358_n13), .IN2(
        DP_OP_342_163_2358_n12), .OUT(C1_DATA4_5) );
  NOR2X1 DP_OP_342_163_2358_U16 ( .IN1(DP_OP_349_170_2358_n58), .IN2(
        DP_OP_342_163_2358_n26), .OUT(DP_OP_342_163_2358_n11) );
  NOR2X1 DP_OP_342_163_2358_U13 ( .IN1(DP_OP_342_163_2358_n26), .IN2(
        DP_OP_342_163_2358_n11), .OUT(DP_OP_342_163_2358_n9) );
  NOR2X1 DP_OP_342_163_2358_U12 ( .IN1(DP_OP_349_170_2358_n58), .IN2(
        DP_OP_342_163_2358_n11), .OUT(DP_OP_342_163_2358_n8) );
  NOR2X1 DP_OP_342_163_2358_U11 ( .IN1(DP_OP_342_163_2358_n9), .IN2(
        DP_OP_342_163_2358_n8), .OUT(C1_DATA4_6) );
  NOR2X1 DP_OP_342_163_2358_U10 ( .IN1(n181), .IN2(DP_OP_342_163_2358_n25), 
        .OUT(DP_OP_342_163_2358_n7) );
  NOR2X1 DP_OP_342_163_2358_U7 ( .IN1(DP_OP_342_163_2358_n25), .IN2(
        DP_OP_342_163_2358_n7), .OUT(DP_OP_342_163_2358_n5) );
  NOR2X1 DP_OP_342_163_2358_U6 ( .IN1(n181), .IN2(DP_OP_342_163_2358_n7), 
        .OUT(DP_OP_342_163_2358_n4) );
  NOR2X1 DP_OP_342_163_2358_U5 ( .IN1(DP_OP_342_163_2358_n5), .IN2(
        DP_OP_342_163_2358_n4), .OUT(C1_DATA4_7) );
  NOR2X1 DP_OP_342_163_2358_U4 ( .IN1(DP_OP_342_163_2358_n24), .IN2(n408), 
        .OUT(DP_OP_342_163_2358_n3) );
  NOR2X1 DP_OP_342_163_2358_U3 ( .IN1(DP_OP_342_163_2358_n24), .IN2(
        DP_OP_342_163_2358_n3), .OUT(DP_OP_342_163_2358_n2) );
  NOR2X1 DP_OP_342_163_2358_U2 ( .IN1(n408), .IN2(DP_OP_342_163_2358_n3), 
        .OUT(DP_OP_342_163_2358_n1) );
  NOR2X1 DP_OP_342_163_2358_U1 ( .IN1(DP_OP_342_163_2358_n2), .IN2(
        DP_OP_342_163_2358_n1), .OUT(C1_DATA4_8) );
  NOR2X1 DP_OP_346_167_2358_U28 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_349_170_2358_n56), .OUT(DP_OP_346_167_2358_n19) );
  NOR2X1 DP_OP_346_167_2358_U25 ( .IN1(DP_OP_349_170_2358_n56), .IN2(
        DP_OP_346_167_2358_n19), .OUT(DP_OP_346_167_2358_n17) );
  NOR2X1 DP_OP_346_167_2358_U24 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_346_167_2358_n19), .OUT(DP_OP_346_167_2358_n16) );
  NOR2X1 DP_OP_346_167_2358_U23 ( .IN1(DP_OP_346_167_2358_n17), .IN2(
        DP_OP_346_167_2358_n16), .OUT(C1_DATA8_4) );
  NOR2X1 DP_OP_346_167_2358_U22 ( .IN1(DP_OP_349_170_2358_n57), .IN2(
        DP_OP_346_167_2358_n23), .OUT(DP_OP_346_167_2358_n15) );
  NOR2X1 DP_OP_346_167_2358_U16 ( .IN1(DP_OP_349_170_2358_n58), .IN2(
        DP_OP_346_167_2358_n22), .OUT(DP_OP_346_167_2358_n11) );
  NOR2X1 DP_OP_346_167_2358_U10 ( .IN1(n181), .IN2(DP_OP_346_167_2358_n21), 
        .OUT(DP_OP_346_167_2358_n7) );
  INVX1 DP_OP_269_159_6943_U91 ( .IN(DP_OP_269_159_6943_n78), .OUT(
        DP_OP_269_159_6943_n76) );
  INVX1 DP_OP_269_159_6943_U6 ( .IN(DP_OP_269_159_6943_n90), .OUT(
        DP_OP_269_159_6943_n29) );
  INVX1 DP_OP_344_165_2358_U33 ( .IN(DP_OP_344_165_2358_n23), .OUT(
        DP_OP_344_165_2358_n32) );
  INVX1 DP_OP_344_165_2358_U9 ( .IN(DP_OP_344_165_2358_n7), .OUT(
        DP_OP_344_165_2358_n28) );
  INVX1 DP_OP_348_169_2358_U21 ( .IN(DP_OP_348_169_2358_n15), .OUT(
        DP_OP_348_169_2358_n30) );
  INVX1 DP_OP_348_169_2358_U15 ( .IN(DP_OP_348_169_2358_n11), .OUT(
        DP_OP_348_169_2358_n29) );
  INVX1 DP_OP_350_171_2358_U27 ( .IN(DP_OP_350_171_2358_n19), .OUT(
        DP_OP_350_171_2358_n27) );
  INVX1 DP_OP_350_171_2358_U21 ( .IN(DP_OP_350_171_2358_n15), .OUT(
        DP_OP_350_171_2358_n26) );
  INVX1 DP_OP_350_171_2358_U15 ( .IN(DP_OP_350_171_2358_n11), .OUT(
        DP_OP_350_171_2358_n25) );
  INVX1 DP_OP_350_171_2358_U9 ( .IN(DP_OP_350_171_2358_n7), .OUT(
        DP_OP_350_171_2358_n24) );
  INVX1 DP_OP_346_167_2358_U27 ( .IN(DP_OP_346_167_2358_n19), .OUT(
        DP_OP_346_167_2358_n23) );
  INVX1 DP_OP_346_167_2358_U21 ( .IN(DP_OP_346_167_2358_n15), .OUT(
        DP_OP_346_167_2358_n22) );
  INVX1 DP_OP_346_167_2358_U15 ( .IN(DP_OP_346_167_2358_n11), .OUT(
        DP_OP_346_167_2358_n21) );
  INVX1 DP_OP_351_172_2358_U15 ( .IN(DP_OP_351_172_2358_n11), .OUT(
        DP_OP_351_172_2358_n33) );
  INVX1 DP_OP_342_163_2358_U15 ( .IN(DP_OP_342_163_2358_n11), .OUT(
        DP_OP_342_163_2358_n25) );
  INVX1 DP_OP_342_163_2358_U9 ( .IN(DP_OP_342_163_2358_n7), .OUT(
        DP_OP_342_163_2358_n24) );
  INVX1 DP_OP_349_170_2358_U15 ( .IN(DP_OP_349_170_2358_n11), .OUT(
        DP_OP_349_170_2358_n33) );
  INVX1 DP_OP_349_170_2358_U9 ( .IN(DP_OP_349_170_2358_n7), .OUT(
        DP_OP_349_170_2358_n32) );
  INVX1 DP_OP_345_166_2358_U21 ( .IN(DP_OP_345_166_2358_n15), .OUT(
        DP_OP_345_166_2358_n34) );
  INVX1 DP_OP_345_166_2358_U15 ( .IN(DP_OP_345_166_2358_n11), .OUT(
        DP_OP_345_166_2358_n33) );
  INVX1 DP_OP_347_168_2358_U27 ( .IN(DP_OP_347_168_2358_n19), .OUT(
        DP_OP_347_168_2358_n35) );
  INVX1 DP_OP_269_159_6943_U27 ( .IN(DP_OP_269_159_6943_n50), .OUT(
        DP_OP_269_159_6943_n48) );
  INVX1 DP_OP_269_159_6943_U28 ( .IN(DP_OP_269_159_6943_n51), .OUT(
        DP_OP_269_159_6943_n49) );
  INVX1 DP_OP_269_159_6943_U17 ( .IN(DP_OP_269_159_6943_n43), .OUT(
        DP_OP_269_159_6943_n79) );
  INVX1 DP_OP_344_165_2358_U27 ( .IN(DP_OP_344_165_2358_n19), .OUT(
        DP_OP_344_165_2358_n31) );
  INVX1 DP_OP_269_159_6943_U82 ( .IN(DP_OP_269_159_6943_n72), .OUT(
        DP_OP_269_159_6943_n85) );
  NAND2X1 DP_OP_351_172_2358_U30 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_351_172_2358_n23), .OUT(DP_OP_351_172_2358_n20) );
  NAND2X1 DP_OP_347_168_2358_U30 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_347_168_2358_n23), .OUT(DP_OP_347_168_2358_n20) );
  NAND2X1 DP_OP_349_170_2358_U30 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_349_170_2358_n23), .OUT(DP_OP_349_170_2358_n20) );
  INVX1 DP_OP_269_159_6943_U79 ( .IN(DP_OP_269_159_6943_n71), .OUT(
        DP_OP_269_159_6943_n70) );
  INVX1 DP_OP_269_159_6943_U63 ( .IN(DP_OP_269_159_6943_n65), .OUT(
        DP_OP_269_159_6943_n83) );
  NAND2X1 DP_OP_351_172_2358_U37 ( .IN1(DP_OP_343_164_2358_n38), .IN2(
        DP_OP_351_172_2358_n27), .OUT(DP_OP_351_172_2358_n25) );
  NAND2X1 DP_OP_351_172_2358_U36 ( .IN1(n394), .IN2(DP_OP_351_172_2358_n27), 
        .OUT(DP_OP_351_172_2358_n24) );
  NAND2X1 DP_OP_343_164_2358_U36 ( .IN1(n394), .IN2(DP_OP_343_164_2358_n27), 
        .OUT(DP_OP_343_164_2358_n24) );
  INVX1 DP_OP_269_159_6943_U52 ( .IN(DP_OP_269_159_6943_n60), .OUT(
        DP_OP_269_159_6943_n82) );
  INVX1 DP_OP_351_172_2358_U33 ( .IN(DP_OP_351_172_2358_n23), .OUT(
        DP_OP_351_172_2358_n36) );
  INVX1 DP_OP_349_170_2358_U33 ( .IN(DP_OP_349_170_2358_n23), .OUT(
        DP_OP_349_170_2358_n36) );
  NANDX2 DP_OP_269_159_6943_U84 ( .IN1(DP_OP_269_159_6943_n103), .IN2(n431), 
        .OUT(DP_OP_269_159_6943_n73) );
  NANDX2 DP_OP_269_159_6943_U74 ( .IN1(DP_OP_269_159_6943_n101), .IN2(
        DP_OP_269_159_6943_n102), .OUT(DP_OP_269_159_6943_n69) );
  NANDX2 DP_OP_269_159_6943_U65 ( .IN1(DP_OP_269_159_6943_n99), .IN2(
        DP_OP_269_159_6943_n100), .OUT(DP_OP_269_159_6943_n66) );
  NANDX2 DP_OP_269_159_6943_U54 ( .IN1(DP_OP_269_159_6943_n97), .IN2(
        DP_OP_269_159_6943_n98), .OUT(DP_OP_269_159_6943_n61) );
  NANDX2 DP_OP_269_159_6943_U32 ( .IN1(DP_OP_269_159_6943_n93), .IN2(
        DP_OP_269_159_6943_n94), .OUT(DP_OP_269_159_6943_n51) );
  INVX4 DP_OP_350_171_2358_U33 ( .IN(DP_OP_350_171_2358_n23), .OUT(
        DP_OP_350_171_2358_n28) );
  INVX4 DP_OP_341_162_2358_U45 ( .IN(DP_OP_345_166_2358_n31), .OUT(
        DP_OP_341_162_2358_n38) );
  INVX4 DP_OP_343_164_2358_U39 ( .IN(DP_OP_343_164_2358_n27), .OUT(
        DP_OP_343_164_2358_n37) );
  INVX4 DP_OP_347_168_2358_U33 ( .IN(DP_OP_347_168_2358_n23), .OUT(
        DP_OP_347_168_2358_n36) );
  NANDX2 DP_OP_349_170_2358_U41 ( .IN1(DP_OP_341_162_2358_n29), .IN2(
        DP_OP_341_162_2358_n28), .OUT(C1_DATA11_1) );
  NANDX2 DP_OP_351_172_2358_U29 ( .IN1(DP_OP_351_172_2358_n21), .IN2(
        DP_OP_351_172_2358_n20), .OUT(C1_DATA13_3) );
  NANDX2 DP_OP_347_168_2358_U29 ( .IN1(DP_OP_347_168_2358_n21), .IN2(
        DP_OP_347_168_2358_n20), .OUT(C1_DATA9_3) );
  NANDX2 DP_OP_349_170_2358_U29 ( .IN1(DP_OP_349_170_2358_n21), .IN2(
        DP_OP_349_170_2358_n20), .OUT(C1_DATA11_3) );
  NANDX2 DP_OP_351_172_2358_U35 ( .IN1(DP_OP_351_172_2358_n25), .IN2(
        DP_OP_351_172_2358_n24), .OUT(C1_DATA13_2) );
  NANDX2 DP_OP_343_164_2358_U35 ( .IN1(DP_OP_343_164_2358_n25), .IN2(
        DP_OP_343_164_2358_n24), .OUT(C1_DATA5_2) );
  NANDX2 DP_OP_351_172_2358_U40 ( .IN1(n394), .IN2(DP_OP_343_164_2358_n38), 
        .OUT(DP_OP_351_172_2358_n27) );
  NANDX2 DP_OP_351_172_2358_U34 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_343_164_2358_n37), .OUT(DP_OP_351_172_2358_n23) );
  INVX1 DP_OP_342_163_2358_U21 ( .IN(DP_OP_342_163_2358_n15), .OUT(
        DP_OP_342_163_2358_n26) );
  NAND2X1 DP_OP_347_168_2358_U31 ( .IN1(DP_OP_347_168_2358_n37), .IN2(
        DP_OP_347_168_2358_n23), .OUT(DP_OP_347_168_2358_n21) );
  NAND2X1 DP_OP_349_170_2358_U31 ( .IN1(DP_OP_341_162_2358_n37), .IN2(
        DP_OP_349_170_2358_n23), .OUT(DP_OP_349_170_2358_n21) );
  NAND2X1 DP_OP_269_159_6943_U19 ( .IN1(DP_OP_269_159_6943_n92), .IN2(
        DP_OP_269_159_6943_n91), .OUT(DP_OP_269_159_6943_n44) );
  NANDX2 DP_OP_349_170_2358_U34 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_341_162_2358_n37), .OUT(DP_OP_349_170_2358_n23) );
  NANDX2 DP_OP_343_164_2358_U40 ( .IN1(n394), .IN2(DP_OP_343_164_2358_n38), 
        .OUT(DP_OP_343_164_2358_n27) );
  NANDX2 DP_OP_347_168_2358_U34 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        DP_OP_347_168_2358_n37), .OUT(DP_OP_347_168_2358_n23) );
  INVX1 DP_OP_269_159_6943_U90 ( .IN(DP_OP_269_159_6943_n77), .OUT(
        DP_OP_269_159_6943_n75) );
  NANDX2 DP_OP_350_171_2358_U34 ( .IN1(DP_OP_349_170_2358_n55), .IN2(
        Final_Exponent_reg[2]), .OUT(DP_OP_350_171_2358_n23) );
  INVX1 DP_OP_344_165_2358_U39 ( .IN(n482), .OUT(DP_OP_344_165_2358_n33) );
  NANDX2 DP_OP_269_159_6943_U12 ( .IN1(DP_OP_269_159_6943_n55), .IN2(
        DP_OP_269_159_6943_n41), .OUT(DP_OP_269_159_6943_n39) );
  NAND2X1 DP_OP_269_159_6943_U62 ( .IN1(DP_OP_269_159_6943_n83), .IN2(
        DP_OP_269_159_6943_n66), .OUT(DP_OP_269_159_6943_n34) );
  NANDX2 DP_OP_351_172_2358_U31 ( .IN1(DP_OP_343_164_2358_n37), .IN2(
        DP_OP_351_172_2358_n23), .OUT(DP_OP_351_172_2358_n21) );
  NANDX2 DP_OP_269_159_6943_U45 ( .IN1(DP_OP_269_159_6943_n95), .IN2(
        DP_OP_269_159_6943_n96), .OUT(DP_OP_269_159_6943_n58) );
  NAND2X1 DP_OP_341_162_2358_U41 ( .IN1(DP_OP_341_162_2358_n29), .IN2(
        DP_OP_341_162_2358_n28), .OUT(C1_DATA3_1) );
  NAND2X1 U3 ( .IN1(DP_OP_344_165_2358_n30), .IN2(DP_OP_349_170_2358_n58), 
        .OUT(n1) );
  NAND2X1 U4 ( .IN1(DP_OP_344_165_2358_n29), .IN2(n1), .OUT(C1_DATA6_6) );
  NAND2X1 U5 ( .IN1(DP_OP_342_163_2358_n28), .IN2(DP_OP_349_170_2358_n56), 
        .OUT(n2) );
  NAND2X1 U6 ( .IN1(n382), .IN2(n2), .OUT(C1_DATA4_4) );
  INVX1 U7 ( .IN(Datain2[9]), .OUT(n3) );
  MUX2X1 U8 ( .IN1(Datain2[9]), .IN2(n3), .S(Datain1[9]), .OUT(
        DP_OP_269_159_6943_n101) );
  OAI21 U9 ( .IN1(n701), .IN2(n4), .IN3(n5), .OUT(n670) );
  INVX1 U10 ( .IN(C1_DATA9_0), .OUT(n4) );
  INVX1 U11 ( .IN(n538), .OUT(n5) );
  INVX1 U12 ( .IN(n408), .OUT(n6) );
  INVX1 U13 ( .IN(DP_OP_346_167_2358_n7), .OUT(n7) );
  AOI22 U14 ( .IN1(DP_OP_346_167_2358_n7), .IN2(n408), .IN3(n6), .IN4(n7), 
        .OUT(C1_DATA8_8) );
  NAND2X1 U15 ( .IN1(N367), .IN2(n842), .OUT(n8) );
  NAND3X1 U16 ( .IN1(n618), .IN2(n617), .IN3(n8), .OUT(n9) );
  AOI21 U17 ( .IN1(n816), .IN2(n181), .IN3(n9), .OUT(n10) );
  NAND2X1 U18 ( .IN1(n785), .IN2(n10), .OUT(n333) );
  AOI21 U19 ( .IN1(DP_OP_349_170_2358_n57), .IN2(DP_OP_340_161_2358_n31), 
        .IN3(DP_OP_340_161_2358_n15), .OUT(n11) );
  AOI22 U20 ( .IN1(n818), .IN2(C1_DATA3_5), .IN3(n817), .IN4(C1_DATA4_5), 
        .OUT(n12) );
  OAI21 U21 ( .IN1(n13), .IN2(n11), .IN3(n12), .OUT(n14) );
  INVX1 U22 ( .IN(n822), .OUT(n13) );
  INVX1 U23 ( .IN(n14), .OUT(n574) );
  INVX1 U24 ( .IN(Datain2[12]), .OUT(n15) );
  MUX2X1 U25 ( .IN1(Datain2[12]), .IN2(n15), .S(Datain1[12]), .OUT(
        DP_OP_269_159_6943_n95) );
  AOI21 U26 ( .IN1(DP_OP_349_170_2358_n56), .IN2(DP_OP_347_168_2358_n36), 
        .IN3(DP_OP_347_168_2358_n19), .OUT(n16) );
  INVX1 U27 ( .IN(n16), .OUT(C1_DATA9_4) );
  INVX1 U28 ( .IN(RSTn_BAR), .OUT(n17) );
  OAI21 U29 ( .IN1(n937), .IN2(n936), .IN3(n935), .OUT(n18) );
  AOI21 U30 ( .IN1(n938), .IN2(Datain2[5]), .IN3(n18), .OUT(n19) );
  OAI21 U31 ( .IN1(n939), .IN2(n958), .IN3(n19), .OUT(n20) );
  AOI22 U32 ( .IN1(Final_Mantissa_reg[5]), .IN2(n959), .IN3(n17), .IN4(n20), 
        .OUT(n21) );
  INVX1 U33 ( .IN(n21), .OUT(n283) );
  OAI21 U34 ( .IN1(DP_OP_341_162_2358_n38), .IN2(n394), .IN3(n468), .OUT(n22)
         );
  INVX1 U35 ( .IN(n22), .OUT(C1_DATA7_2) );
  NAND3X1 U36 ( .IN1(Multi_dataout[14]), .IN2(n803), .IN3(n735), .OUT(n910) );
  INVX1 U37 ( .IN(n408), .OUT(n23) );
  MUX2X1 U38 ( .IN1(n23), .IN2(n408), .S(DP_OP_339_160_2358_n32), .OUT(
        C1_DATA1_8) );
  INVX1 U39 ( .IN(n408), .OUT(n24) );
  MUX2X1 U40 ( .IN1(n24), .IN2(n408), .S(DP_OP_344_165_2358_n28), .OUT(
        C1_DATA6_8) );
  NAND2X1 U41 ( .IN1(DP_OP_269_159_6943_n61), .IN2(DP_OP_269_159_6943_n82), 
        .OUT(n25) );
  AOI22 U42 ( .IN1(Datain1[11]), .IN2(n916), .IN3(Datain2[11]), .IN4(n957), 
        .OUT(n26) );
  INVX1 U43 ( .IN(DP_OP_269_159_6943_n62), .OUT(n27) );
  MUX2X1 U44 ( .IN1(n27), .IN2(DP_OP_269_159_6943_n62), .S(n25), .OUT(n28) );
  OAI21 U45 ( .IN1(n619), .IN2(n28), .IN3(n26), .OUT(n598) );
  NAND2X1 U46 ( .IN1(DP_OP_340_161_2358_n32), .IN2(DP_OP_349_170_2358_n56), 
        .OUT(n29) );
  NAND2X1 U47 ( .IN1(DP_OP_340_161_2358_n31), .IN2(n29), .OUT(C1_DATA2_4) );
  NAND2X1 U48 ( .IN1(DP_OP_347_168_2358_n38), .IN2(n394), .OUT(n30) );
  NAND2X1 U49 ( .IN1(DP_OP_347_168_2358_n37), .IN2(n30), .OUT(C1_DATA9_2) );
  AOI22 U50 ( .IN1(n412), .IN2(Datain1[8]), .IN3(n423), .IN4(Datain2[8]), 
        .OUT(n31) );
  INVX1 U51 ( .IN(n31), .OUT(DP_OP_269_159_6943_n103) );
  INVX1 U52 ( .IN(n956), .OUT(n32) );
  AOI22 U53 ( .IN1(n954), .IN2(n955), .IN3(Datain1[6]), .IN4(n32), .OUT(n33)
         );
  NAND2X1 U54 ( .IN1(n409), .IN2(Multi_dataout[14]), .OUT(n34) );
  OAI21 U55 ( .IN1(n958), .IN2(n34), .IN3(n33), .OUT(n35) );
  AOI21 U56 ( .IN1(n957), .IN2(Datain2[6]), .IN3(n35), .OUT(n36) );
  NAND2X1 U57 ( .IN1(n959), .IN2(Final_Mantissa_reg[6]), .OUT(n37) );
  NAND2X1 U58 ( .IN1(n36), .IN2(n37), .OUT(n345) );
  INVX1 U59 ( .IN(DP_OP_349_170_2358_n58), .OUT(n38) );
  NAND2X1 U60 ( .IN1(DP_OP_343_164_2358_n15), .IN2(n38), .OUT(n162) );
  NAND3X1 U61 ( .IN1(Final_Mantissa_reg[0]), .IN2(Final_Mantissa_reg[1]), 
        .IN3(G_reg), .OUT(n39) );
  INVX1 U62 ( .IN(n39), .OUT(n890) );
  OAI21 U63 ( .IN1(n404), .IN2(n394), .IN3(n482), .OUT(n40) );
  INVX1 U64 ( .IN(n40), .OUT(C1_DATA6_2) );
  NAND2X1 U65 ( .IN1(DP_OP_269_159_6943_n44), .IN2(DP_OP_269_159_6943_n79), 
        .OUT(n41) );
  INVX1 U66 ( .IN(n41), .OUT(n42) );
  AOI21 U67 ( .IN1(DP_OP_269_159_6943_n56), .IN2(DP_OP_269_159_6943_n48), 
        .IN3(DP_OP_269_159_6943_n49), .OUT(n43) );
  OAI21 U68 ( .IN1(DP_OP_269_159_6943_n62), .IN2(DP_OP_269_159_6943_n46), 
        .IN3(n43), .OUT(n44) );
  MUX2X1 U69 ( .IN1(n42), .IN2(n41), .S(n44), .OUT(N367) );
  INVX1 U70 ( .IN(DP_OP_347_168_2358_n7), .OUT(n45) );
  MUX2X1 U71 ( .IN1(DP_OP_347_168_2358_n7), .IN2(n45), .S(n408), .OUT(
        C1_DATA9_8) );
  INVX1 U72 ( .IN(DP_OP_348_169_2358_n7), .OUT(n46) );
  MUX2X1 U73 ( .IN1(DP_OP_348_169_2358_n7), .IN2(n46), .S(n408), .OUT(
        C1_DATA10_8) );
  NAND3X1 U74 ( .IN1(n180), .IN2(n186), .IN3(n192), .OUT(n445) );
  AOI21 U75 ( .IN1(Datain1[14]), .IN2(Datain2[14]), .IN3(
        DP_OP_269_159_6943_n90), .OUT(n47) );
  INVX1 U76 ( .IN(n47), .OUT(DP_OP_269_159_6943_n91) );
  INVX1 U77 ( .IN(DP_OP_349_170_2358_n58), .OUT(n48) );
  OAI21 U78 ( .IN1(DP_OP_343_164_2358_n15), .IN2(n48), .IN3(n162), .OUT(
        C1_DATA5_6) );
  AOI21 U79 ( .IN1(DP_OP_349_170_2358_n58), .IN2(DP_OP_350_171_2358_n26), 
        .IN3(DP_OP_350_171_2358_n11), .OUT(n49) );
  INVX1 U80 ( .IN(n49), .OUT(C1_DATA12_6) );
  NAND3X1 U81 ( .IN1(n334), .IN2(n540), .IN3(n863), .OUT(n50) );
  NOR2X1 U82 ( .IN1(n285), .IN2(n50), .OUT(n542) );
  AOI21 U83 ( .IN1(n181), .IN2(DP_OP_345_166_2358_n33), .IN3(
        DP_OP_345_166_2358_n7), .OUT(n51) );
  INVX1 U84 ( .IN(n51), .OUT(C1_DATA7_7) );
  AOI21 U85 ( .IN1(n181), .IN2(DP_OP_351_172_2358_n33), .IN3(
        DP_OP_351_172_2358_n7), .OUT(n52) );
  INVX1 U86 ( .IN(n52), .OUT(C1_DATA13_7) );
  AOI21 U87 ( .IN1(C1_DATA8_0), .IN2(n404), .IN3(DP_OP_347_168_2358_n31), 
        .OUT(n53) );
  INVX1 U88 ( .IN(n53), .OUT(n54) );
  AOI22 U89 ( .IN1(n826), .IN2(n54), .IN3(C1_DATA11_1), .IN4(n827), .OUT(n563)
         );
  AOI21 U90 ( .IN1(Exc_value[2]), .IN2(n193), .IN3(n456), .OUT(n55) );
  INVX1 U91 ( .IN(n55), .OUT(n549) );
  NAND2X1 U92 ( .IN1(DP_OP_269_159_6943_n51), .IN2(DP_OP_269_159_6943_n48), 
        .OUT(n56) );
  INVX1 U93 ( .IN(n56), .OUT(n57) );
  INVX1 U94 ( .IN(DP_OP_269_159_6943_n62), .OUT(n58) );
  AOI21 U95 ( .IN1(DP_OP_269_159_6943_n55), .IN2(n58), .IN3(
        DP_OP_269_159_6943_n56), .OUT(n60) );
  MUX2X1 U96 ( .IN1(n56), .IN2(n57), .S(n60), .OUT(N366) );
  INVX1 U97 ( .IN(n277), .OUT(n61) );
  NAND3X1 U98 ( .IN1(Multi_dataout[0]), .IN2(n271), .IN3(n61), .OUT(n62) );
  NAND3X1 U99 ( .IN1(n875), .IN2(n876), .IN3(n62), .OUT(n877) );
  AOI22 U100 ( .IN1(Datain1[10]), .IN2(n916), .IN3(Datain2[10]), .IN4(n957), 
        .OUT(n63) );
  NAND3X1 U101 ( .IN1(n650), .IN2(n781), .IN3(n649), .OUT(n64) );
  NAND2X1 U102 ( .IN1(n63), .IN2(n64), .OUT(n65) );
  INVX1 U103 ( .IN(DP_OP_269_159_6943_n67), .OUT(n66) );
  MUX2X1 U104 ( .IN1(n66), .IN2(DP_OP_269_159_6943_n67), .S(
        DP_OP_269_159_6943_n34), .OUT(n67) );
  AOI21 U105 ( .IN1(n67), .IN2(n842), .IN3(n65), .OUT(n651) );
  NAND2X1 U106 ( .IN1(Datain2[13]), .IN2(Datain1[13]), .OUT(n68) );
  INVX1 U107 ( .IN(n68), .OUT(DP_OP_269_159_6943_n92) );
  NAND3X1 U108 ( .IN1(n328), .IN2(n712), .IN3(n268), .OUT(n373) );
  NAND2X1 U109 ( .IN1(DP_OP_341_162_2358_n37), .IN2(DP_OP_349_170_2358_n55), 
        .OUT(n69) );
  OAI21 U110 ( .IN1(DP_OP_341_162_2358_n23), .IN2(n70), .IN3(n818), .OUT(n639)
         );
  INVX1 U111 ( .IN(n69), .OUT(n70) );
  MUX2X1 U112 ( .IN1(Datain1[10]), .IN2(n427), .S(Datain2[10]), .OUT(
        DP_OP_269_159_6943_n99) );
  AOI21 U113 ( .IN1(DP_OP_349_170_2358_n58), .IN2(DP_OP_347_168_2358_n34), 
        .IN3(DP_OP_347_168_2358_n11), .OUT(n71) );
  INVX1 U114 ( .IN(n71), .OUT(C1_DATA9_6) );
  AOI21 U115 ( .IN1(DP_OP_349_170_2358_n58), .IN2(DP_OP_346_167_2358_n22), 
        .IN3(DP_OP_346_167_2358_n11), .OUT(n72) );
  INVX1 U116 ( .IN(n72), .OUT(C1_DATA8_6) );
  NAND3X1 U117 ( .IN1(DP_OP_349_170_2358_n57), .IN2(n599), .IN3(
        DP_OP_349_170_2358_n56), .OUT(n603) );
  NAND2X1 U118 ( .IN1(DP_OP_343_164_2358_n36), .IN2(DP_OP_349_170_2358_n56), 
        .OUT(n73) );
  NAND2X1 U119 ( .IN1(n398), .IN2(n73), .OUT(C1_DATA5_4) );
  MUX2X1 U120 ( .IN1(Datain1[11]), .IN2(n426), .S(Datain2[11]), .OUT(
        DP_OP_269_159_6943_n97) );
  NAND3X1 U121 ( .IN1(Final_Mantissa_reg[4]), .IN2(n924), .IN3(
        Final_Mantissa_reg[5]), .OUT(n953) );
  AOI21 U122 ( .IN1(n181), .IN2(DP_OP_349_170_2358_n33), .IN3(
        DP_OP_349_170_2358_n7), .OUT(n74) );
  INVX1 U123 ( .IN(n74), .OUT(C1_DATA11_7) );
  AOI21 U124 ( .IN1(n181), .IN2(DP_OP_350_171_2358_n25), .IN3(
        DP_OP_350_171_2358_n7), .OUT(n75) );
  INVX1 U125 ( .IN(n75), .OUT(C1_DATA12_7) );
  OAI21 U126 ( .IN1(n544), .IN2(n242), .IN3(n409), .OUT(n76) );
  NAND3X1 U127 ( .IN1(n724), .IN2(n718), .IN3(n542), .OUT(n77) );
  NOR2X1 U128 ( .IN1(n544), .IN2(Multi_dataout[14]), .OUT(n78) );
  AOI21 U129 ( .IN1(n78), .IN2(n77), .IN3(n76), .OUT(n79) );
  INVX1 U130 ( .IN(n79), .OUT(n239) );
  INVX1 U131 ( .IN(RSOP_340_C1_Z_0), .OUT(n80) );
  NAND2X1 U132 ( .IN1(DP_OP_269_159_6943_n78), .IN2(DP_OP_269_159_6943_n75), 
        .OUT(n81) );
  MUX2X1 U133 ( .IN1(n80), .IN2(RSOP_340_C1_Z_0), .S(n81), .OUT(N360) );
  INVX1 U134 ( .IN(DP_OP_345_166_2358_n7), .OUT(n82) );
  MUX2X1 U135 ( .IN1(DP_OP_345_166_2358_n7), .IN2(n82), .S(n408), .OUT(
        C1_DATA7_8) );
  INVX1 U136 ( .IN(DP_OP_351_172_2358_n7), .OUT(n83) );
  MUX2X1 U137 ( .IN1(DP_OP_351_172_2358_n7), .IN2(n83), .S(n408), .OUT(
        C1_DATA13_8) );
  INVX1 U138 ( .IN(n960), .OUT(n84) );
  NOR2X1 U139 ( .IN1(n296), .IN2(n84), .OUT(n330) );
  AOI22 U140 ( .IN1(Datain1[9]), .IN2(n916), .IN3(Datain2[9]), .IN4(n957), 
        .OUT(n85) );
  INVX1 U141 ( .IN(DP_OP_269_159_6943_n68), .OUT(n86) );
  NAND2X1 U142 ( .IN1(DP_OP_269_159_6943_n69), .IN2(n86), .OUT(n87) );
  INVX1 U143 ( .IN(DP_OP_269_159_6943_n70), .OUT(n88) );
  MUX2X1 U144 ( .IN1(n88), .IN2(DP_OP_269_159_6943_n70), .S(n87), .OUT(n90) );
  OAI21 U145 ( .IN1(n619), .IN2(n90), .IN3(n85), .OUT(n633) );
  INVX1 U146 ( .IN(n549), .OUT(n91) );
  INVX1 U147 ( .IN(n551), .OUT(n92) );
  NAND3X1 U148 ( .IN1(n550), .IN2(n91), .IN3(n92), .OUT(n850) );
  NAND3X1 U149 ( .IN1(n676), .IN2(n720), .IN3(n675), .OUT(n273) );
  AOI21 U150 ( .IN1(DP_OP_349_170_2358_n58), .IN2(DP_OP_341_162_2358_n34), 
        .IN3(DP_OP_341_162_2358_n11), .OUT(n93) );
  INVX1 U151 ( .IN(n93), .OUT(C1_DATA3_6) );
  INVX1 U152 ( .IN(n491), .OUT(n94) );
  AOI21 U153 ( .IN1(n462), .IN2(n499), .IN3(n94), .OUT(n369) );
  AOI21 U154 ( .IN1(DP_OP_349_170_2358_n58), .IN2(DP_OP_345_166_2358_n34), 
        .IN3(DP_OP_345_166_2358_n11), .OUT(n95) );
  INVX1 U155 ( .IN(n95), .OUT(C1_DATA7_6) );
  AOI21 U156 ( .IN1(DP_OP_349_170_2358_n58), .IN2(DP_OP_348_169_2358_n30), 
        .IN3(DP_OP_348_169_2358_n11), .OUT(n98) );
  INVX1 U157 ( .IN(n98), .OUT(C1_DATA10_6) );
  AOI21 U158 ( .IN1(n115), .IN2(n131), .IN3(DP_OP_350_171_2358_n13), .OUT(n132) );
  AOI21 U159 ( .IN1(DP_OP_349_170_2358_n57), .IN2(DP_OP_346_167_2358_n23), 
        .IN3(DP_OP_346_167_2358_n15), .OUT(n133) );
  INVX1 U160 ( .IN(n133), .OUT(n134) );
  AOI22 U161 ( .IN1(n834), .IN2(n132), .IN3(n833), .IN4(n134), .OUT(n576) );
  INVX1 U162 ( .IN(DP_OP_349_170_2358_n57), .OUT(n115) );
  INVX1 U163 ( .IN(DP_OP_350_171_2358_n15), .OUT(n131) );
  NAND3X1 U164 ( .IN1(Final_Mantissa_reg[3]), .IN2(n890), .IN3(
        Final_Mantissa_reg[2]), .OUT(n933) );
  OAI21 U165 ( .IN1(n394), .IN2(DP_OP_349_170_2358_n55), .IN3(
        DP_OP_350_171_2358_n23), .OUT(n135) );
  INVX1 U166 ( .IN(n135), .OUT(C1_DATA12_3) );
  NAND3X1 U167 ( .IN1(n178), .IN2(DP_OP_339_160_2358_n15), .IN3(n184), .OUT(
        DP_OP_339_160_2358_n32) );
  AOI21 U168 ( .IN1(n181), .IN2(DP_OP_347_168_2358_n33), .IN3(
        DP_OP_347_168_2358_n7), .OUT(n136) );
  INVX1 U169 ( .IN(n136), .OUT(C1_DATA9_7) );
  AOI21 U170 ( .IN1(n181), .IN2(DP_OP_346_167_2358_n21), .IN3(
        DP_OP_346_167_2358_n7), .OUT(n137) );
  INVX1 U171 ( .IN(n137), .OUT(C1_DATA8_7) );
  AOI21 U172 ( .IN1(DP_OP_349_170_2358_n56), .IN2(DP_OP_349_170_2358_n36), 
        .IN3(DP_OP_349_170_2358_n19), .OUT(n138) );
  AOI21 U173 ( .IN1(DP_OP_349_170_2358_n56), .IN2(DP_OP_339_160_2358_n36), 
        .IN3(DP_OP_339_160_2358_n19), .OUT(n139) );
  INVX1 U174 ( .IN(n139), .OUT(n140) );
  NOR2X1 U175 ( .IN1(DP_OP_341_162_2358_n17), .IN2(DP_OP_341_162_2358_n16), 
        .OUT(n141) );
  AOI22 U176 ( .IN1(n820), .IN2(n140), .IN3(n818), .IN4(n141), .OUT(n142) );
  OAI21 U177 ( .IN1(n728), .IN2(n138), .IN3(n142), .OUT(n594) );
  AOI21 U178 ( .IN1(DP_OP_349_170_2358_n55), .IN2(DP_OP_344_165_2358_n33), 
        .IN3(DP_OP_344_165_2358_n23), .OUT(n143) );
  INVX1 U179 ( .IN(n143), .OUT(n144) );
  OAI21 U180 ( .IN1(DP_OP_349_170_2358_n55), .IN2(n174), .IN3(
        DP_OP_348_169_2358_n23), .OUT(n145) );
  INVX1 U181 ( .IN(n145), .OUT(n146) );
  AOI22 U182 ( .IN1(n832), .IN2(n144), .IN3(n831), .IN4(n146), .OUT(n646) );
  NAND3X1 U183 ( .IN1(n181), .IN2(n782), .IN3(DP_OP_349_170_2358_n58), .OUT(
        n605) );
  NOR2X1 U184 ( .IN1(DP_OP_269_159_6943_n57), .IN2(n147), .OUT(n148) );
  INVX1 U185 ( .IN(n148), .OUT(n149) );
  OAI21 U186 ( .IN1(DP_OP_269_159_6943_n62), .IN2(DP_OP_269_159_6943_n60), 
        .IN3(DP_OP_269_159_6943_n61), .OUT(n150) );
  MUX2X1 U187 ( .IN1(n148), .IN2(n149), .S(n150), .OUT(N365) );
  INVX1 U188 ( .IN(DP_OP_269_159_6943_n58), .OUT(n147) );
  INVX1 U189 ( .IN(DP_OP_269_159_6943_n74), .OUT(n151) );
  NAND2X1 U190 ( .IN1(DP_OP_269_159_6943_n73), .IN2(DP_OP_269_159_6943_n85), 
        .OUT(n152) );
  MUX2X1 U191 ( .IN1(DP_OP_269_159_6943_n74), .IN2(n151), .S(n152), .OUT(n153)
         );
  AOI22 U192 ( .IN1(Datain2[8]), .IN2(n957), .IN3(Datain1[8]), .IN4(n916), 
        .OUT(n154) );
  NAND3X1 U193 ( .IN1(C1_DATA8_0), .IN2(n781), .IN3(DP_OP_345_166_2358_n31), 
        .OUT(n155) );
  NAND2X1 U194 ( .IN1(n154), .IN2(n155), .OUT(n156) );
  AOI21 U195 ( .IN1(n842), .IN2(n153), .IN3(n156), .OUT(n565) );
  INVX1 U196 ( .IN(DP_OP_269_159_6943_n3), .OUT(n157) );
  OAI21 U197 ( .IN1(DP_OP_269_159_6943_n29), .IN2(DP_OP_269_159_6943_n4), 
        .IN3(n157), .OUT(n788) );
  INVX1 U198 ( .IN(n705), .OUT(n484) );
  NANDX2 U199 ( .IN1(n471), .IN2(Multi_dataout[11]), .OUT(n349) );
  NAND2X1 U200 ( .IN1(DP_OP_345_166_2358_n31), .IN2(n663), .OUT(n498) );
  BUF4X U201 ( .IN(n478), .OUT(n158) );
  INVX4 U202 ( .IN(n471), .OUT(n159) );
  INVX4 U203 ( .IN(DP_OP_341_162_2358_n27), .OUT(DP_OP_341_162_2358_n37) );
  INVX1 U204 ( .IN(n219), .OUT(n160) );
  INVX4 U205 ( .IN(n219), .OUT(n278) );
  NANDX2 U206 ( .IN1(n668), .IN2(n667), .OUT(n161) );
  NAND2X1 U207 ( .IN1(n668), .IN2(n667), .OUT(n719) );
  INVX1 U208 ( .IN(n251), .OUT(n163) );
  INVX8 U209 ( .IN(n295), .OUT(n168) );
  NANDX2 U210 ( .IN1(n265), .IN2(n260), .OUT(n164) );
  INVX1 U211 ( .IN(n664), .OUT(n822) );
  NAND2X1 U212 ( .IN1(n681), .IN2(n664), .OUT(n665) );
  NAND2X1 U213 ( .IN1(n496), .IN2(n501), .OUT(n681) );
  INVX4 U214 ( .IN(DP_OP_351_172_2358_n31), .OUT(DP_OP_343_164_2358_n38) );
  INVX4 U215 ( .IN(n407), .OUT(DP_OP_349_170_2358_n55) );
  NAND2X1 U216 ( .IN1(n705), .IN2(n863), .OUT(n312) );
  NANDX2 U217 ( .IN1(Multi_dataout[10]), .IN2(n470), .OUT(n208) );
  NAND2X1 U218 ( .IN1(Multi_dataout[8]), .IN2(n163), .OUT(n233) );
  NANDX2 U219 ( .IN1(n175), .IN2(DP_OP_341_162_2358_n23), .OUT(n167) );
  INVX1 U220 ( .IN(n167), .OUT(DP_OP_341_162_2358_n19) );
  INVX4 U221 ( .IN(n251), .OUT(n170) );
  INVX1 U222 ( .IN(n732), .OUT(n835) );
  BUF8X U223 ( .IN(Multi_dataout[5]), .OUT(n391) );
  INVX1 U224 ( .IN(n681), .OUT(n497) );
  INVX1 U225 ( .IN(n208), .OUT(n496) );
  NANDX2 U226 ( .IN1(n263), .IN2(n724), .OUT(n262) );
  NANDX2 U227 ( .IN1(n679), .IN2(n680), .OUT(n261) );
  NAND2X1 U228 ( .IN1(n502), .IN2(n501), .OUT(n533) );
  INVX1 U229 ( .IN(n317), .OUT(n826) );
  NAND2X1 U230 ( .IN1(n729), .IN2(n317), .OUT(n861) );
  INVX1 U231 ( .IN(n728), .OUT(n825) );
  NAND2X1 U232 ( .IN1(n744), .IN2(n743), .OUT(n948) );
  NAND2X1 U233 ( .IN1(Multi_dataout[10]), .IN2(n163), .OUT(n210) );
  BUF8X U234 ( .IN(Multi_dataout[7]), .OUT(n403) );
  NAND2X1 U235 ( .IN1(n288), .IN2(n541), .OUT(n285) );
  NAND2X1 U236 ( .IN1(n479), .IN2(n502), .OUT(n313) );
  NAND2X1 U237 ( .IN1(n391), .IN2(n492), .OUT(n541) );
  NAND2X1 U238 ( .IN1(n308), .IN2(n492), .OUT(n720) );
  BUF4X U239 ( .IN(DP_OP_351_172_2358_n31), .OUT(n169) );
  NANDX2 U240 ( .IN1(n946), .IN2(n925), .OUT(n254) );
  NAND2X1 U241 ( .IN1(n588), .IN2(n587), .OUT(n589) );
  NANDX2 U242 ( .IN1(n311), .IN2(n674), .OUT(n310) );
  NANDX2 U243 ( .IN1(n801), .IN2(n758), .OUT(n799) );
  NANDX2 U244 ( .IN1(n1012), .IN2(n1015), .OUT(n738) );
  NANDX2 U245 ( .IN1(DP_OP_349_170_2358_n55), .IN2(DP_OP_341_162_2358_n38), 
        .OUT(n494) );
  NAND2X1 U246 ( .IN1(n1037), .IN2(n409), .OUT(n1038) );
  INVX1 U247 ( .IN(n992), .OUT(Exc[1]) );
  NANDX2 U248 ( .IN1(n434), .IN2(Data_valid), .OUT(n1043) );
  NAND2X1 U249 ( .IN1(n202), .IN2(Dataout_valid), .OUT(n992) );
  NANDX2 U250 ( .IN1(n303), .IN2(n302), .OUT(n690) );
  NANDX2 U251 ( .IN1(n254), .IN2(n253), .OUT(n252) );
  INVX1 U252 ( .IN(n900), .OUT(n298) );
  INVX1 U253 ( .IN(n256), .OUT(n255) );
  NANDX2 U254 ( .IN1(Multi_dataout[8]), .IN2(n271), .OUT(n246) );
  INVX4 U255 ( .IN(n740), .OUT(n171) );
  NAND2X1 U256 ( .IN1(Multi_dataout[11]), .IN2(n960), .OUT(n926) );
  INVX4 U257 ( .IN(n301), .OUT(n172) );
  INVX1 U258 ( .IN(n284), .OUT(n281) );
  NANDX2 U259 ( .IN1(n739), .IN2(n947), .OUT(n746) );
  NANDX2 U260 ( .IN1(DP_OP_349_170_2358_n57), .IN2(n238), .OUT(n585) );
  NANDX2 U261 ( .IN1(n951), .IN2(n950), .OUT(n964) );
  NANDX2 U262 ( .IN1(n779), .IN2(n778), .OUT(n780) );
  NANDX2 U263 ( .IN1(n240), .IN2(n239), .OUT(n238) );
  NANDX2 U264 ( .IN1(n793), .IN2(n792), .OUT(n794) );
  INVX4 U265 ( .IN(n264), .OUT(n263) );
  NANDX2 U266 ( .IN1(n857), .IN2(n856), .OUT(n858) );
  INVX4 U267 ( .IN(n711), .OUT(n827) );
  NANDX2 U268 ( .IN1(n493), .IN2(n660), .OUT(n729) );
  NANDX2 U269 ( .IN1(n395), .IN2(n922), .OUT(n875) );
  NAND2X1 U270 ( .IN1(C1_DATA3_1), .IN2(n818), .OUT(n555) );
  NANDX2 U271 ( .IN1(C1_DATA5_4), .IN2(n821), .OUT(n591) );
  NAND2X1 U272 ( .IN1(C1_DATA3_2), .IN2(n818), .OUT(n621) );
  INVX1 U273 ( .IN(n736), .OUT(n737) );
  INVX1 U274 ( .IN(DP_OP_339_160_2358_n32), .OUT(DP_OP_339_160_2358_n7) );
  NANDX2 U275 ( .IN1(n505), .IN2(n662), .OUT(n713) );
  INVX1 U276 ( .IN(n539), .OUT(n540) );
  INVX1 U277 ( .IN(n1069), .OUT(n108) );
  INVX1 U278 ( .IN(n1068), .OUT(n109) );
  INVX1 U279 ( .IN(n1066), .OUT(n111) );
  INVX1 U280 ( .IN(n1067), .OUT(n110) );
  INVX1 U281 ( .IN(n522), .OUT(n523) );
  INVX1 U282 ( .IN(n1065), .OUT(n112) );
  INVX1 U283 ( .IN(n1070), .OUT(n107) );
  INVX1 U284 ( .IN(n1072), .OUT(n105) );
  INVX1 U285 ( .IN(n1073), .OUT(n104) );
  INVX1 U286 ( .IN(n1071), .OUT(n106) );
  INVX1 U287 ( .IN(n1074), .OUT(n103) );
  INVX1 U288 ( .IN(n1075), .OUT(n102) );
  INVX1 U289 ( .IN(n1076), .OUT(n101) );
  INVX1 U290 ( .IN(n1077), .OUT(n100) );
  INVX1 U291 ( .IN(n1080), .OUT(n99) );
  INVX1 U292 ( .IN(n1063), .OUT(n114) );
  INVX1 U293 ( .IN(n1064), .OUT(n113) );
  NANDX2 U294 ( .IN1(T_reg), .IN2(n749), .OUT(n355) );
  INVX1 U295 ( .IN(n813), .OUT(n814) );
  NANDX2 U296 ( .IN1(Multi_dataout[15]), .IN2(n803), .OUT(n805) );
  NANDX2 U297 ( .IN1(Final_Mantissa_reg[6]), .IN2(n451), .OUT(n954) );
  INVX1 U298 ( .IN(n1056), .OUT(n119) );
  INVX1 U299 ( .IN(n1055), .OUT(n120) );
  INVX1 U300 ( .IN(n1054), .OUT(n121) );
  INVX1 U301 ( .IN(n1053), .OUT(n122) );
  INVX1 U302 ( .IN(n972), .OUT(n123) );
  INVX1 U303 ( .IN(n1046), .OUT(n130) );
  INVX1 U304 ( .IN(n1047), .OUT(n129) );
  INVX1 U305 ( .IN(n1048), .OUT(n128) );
  INVX1 U306 ( .IN(n1049), .OUT(n127) );
  INVX1 U307 ( .IN(n1050), .OUT(n126) );
  INVX1 U308 ( .IN(n1052), .OUT(n124) );
  INVX1 U309 ( .IN(n1051), .OUT(n125) );
  INVX1 U310 ( .IN(n1060), .OUT(n116) );
  NAND2X1 U311 ( .IN1(n409), .IN2(n938), .OUT(n520) );
  INVX1 U312 ( .IN(n1057), .OUT(n118) );
  INVX1 U313 ( .IN(DP_OP_343_164_2358_n36), .OUT(n176) );
  INVX1 U314 ( .IN(n1058), .OUT(n117) );
  INVX4 U315 ( .IN(n399), .OUT(n395) );
  INVX1 U316 ( .IN(n709), .OUT(n489) );
  NANDX2 U317 ( .IN1(n468), .IN2(n661), .OUT(n475) );
  INVX1 U318 ( .IN(n300), .OUT(n299) );
  NANDX2 U319 ( .IN1(n493), .IN2(n485), .OUT(n659) );
  INVX1 U320 ( .IN(n1003), .OUT(Dataout[9]) );
  NANDX2 U321 ( .IN1(n207), .IN2(n1043), .OUT(n1044) );
  INVX1 U322 ( .IN(n907), .OUT(n909) );
  INVX4 U323 ( .IN(n880), .OUT(n241) );
  INVX1 U324 ( .IN(n991), .OUT(Exc[0]) );
  INVX1 U325 ( .IN(n994), .OUT(Dataout[0]) );
  INVX1 U326 ( .IN(n995), .OUT(Dataout[1]) );
  INVX1 U327 ( .IN(n996), .OUT(Dataout[2]) );
  INVX1 U328 ( .IN(n997), .OUT(Dataout[3]) );
  INVX1 U329 ( .IN(n1008), .OUT(Dataout[14]) );
  INVX1 U330 ( .IN(n1004), .OUT(Dataout[10]) );
  INVX1 U331 ( .IN(n993), .OUT(Exc[2]) );
  INVX1 U332 ( .IN(n1002), .OUT(Dataout[8]) );
  INVX1 U333 ( .IN(n1005), .OUT(Dataout[11]) );
  INVX1 U334 ( .IN(n1006), .OUT(Dataout[12]) );
  INVX1 U335 ( .IN(n1001), .OUT(Dataout[7]) );
  INVX1 U336 ( .IN(n1000), .OUT(Dataout[6]) );
  INVX1 U337 ( .IN(n1007), .OUT(Dataout[13]) );
  INVX1 U338 ( .IN(n999), .OUT(Dataout[5]) );
  INVX1 U339 ( .IN(n998), .OUT(Dataout[4]) );
  NANDX2 U340 ( .IN1(n409), .IN2(n527), .OUT(n880) );
  NAND2X1 U341 ( .IN1(n809), .IN2(n439), .OUT(n754) );
  INVX1 U342 ( .IN(n952), .OUT(n904) );
  NANDX2 U343 ( .IN1(Exc_Ack), .IN2(n987), .OUT(n551) );
  INVX1 U344 ( .IN(n428), .OUT(n429) );
  INVX1 U345 ( .IN(n812), .OUT(n517) );
  INVX1 U346 ( .IN(DP_OP_340_161_2358_n27), .OUT(n174) );
  INVX1 U347 ( .IN(n418), .OUT(n419) );
  NANDX2 U348 ( .IN1(n191), .IN2(n432), .OUT(n1034) );
  INVX1 U349 ( .IN(n990), .OUT(n1010) );
  NANDX2 U350 ( .IN1(StateMC_0_), .IN2(n1014), .OUT(n1040) );
  INVX1 U351 ( .IN(n966), .OUT(n1032) );
  NANDX2 U352 ( .IN1(n203), .IN2(n1016), .OUT(n550) );
  INVX4 U353 ( .IN(C1_DATA8_0), .OUT(C1_DATA9_0) );
  NANDX2 U354 ( .IN1(n179), .IN2(n192), .OUT(n1035) );
  NANDX2 U355 ( .IN1(n188), .IN2(n201), .OUT(n966) );
  INVX4 U356 ( .IN(DP_OP_349_170_2358_n56), .OUT(n175) );
  NANDX2 U357 ( .IN1(n186), .IN2(n437), .OUT(n990) );
  NANDX2 U358 ( .IN1(Multi_dataout[2]), .IN2(n347), .OUT(n674) );
  NAND2X1 U359 ( .IN1(n184), .IN2(DP_OP_339_160_2358_n15), .OUT(
        DP_OP_339_160_2358_n33) );
  NAND2X1 U360 ( .IN1(DP_OP_341_162_2358_n11), .IN2(n178), .OUT(n177) );
  INVX1 U361 ( .IN(n177), .OUT(DP_OP_341_162_2358_n7) );
  BUF4X U362 ( .IN(Final_Exponent_reg[7]), .OUT(n181) );
  INVX1 U363 ( .IN(n671), .OUT(n669) );
  NOR2X1 U364 ( .IN1(n313), .IN2(n314), .OUT(n182) );
  NANDX2 U365 ( .IN1(n501), .IN2(n472), .OUT(n314) );
  INVX1 U366 ( .IN(n725), .OUT(n226) );
  NANDX2 U367 ( .IN1(n725), .IN2(n710), .OUT(n264) );
  INVX1 U368 ( .IN(n312), .OUT(n276) );
  NANDX2 U369 ( .IN1(n946), .IN2(n294), .OUT(n214) );
  NANDX2 U370 ( .IN1(n231), .IN2(n229), .OUT(n688) );
  NAND2X1 U371 ( .IN1(n166), .IN2(DP_OP_347_168_2358_n31), .OUT(
        DP_OP_347_168_2358_n37) );
  NANDX2 U372 ( .IN1(DP_OP_349_170_2358_n55), .IN2(n174), .OUT(
        DP_OP_348_169_2358_n23) );
  NANDX2 U373 ( .IN1(n929), .IN2(n928), .OUT(n689) );
  NANDX2 U374 ( .IN1(n214), .IN2(n211), .OUT(n374) );
  INVX4 U375 ( .IN(n805), .OUT(n848) );
  INVX4 U376 ( .IN(n1034), .OUT(n801) );
  INVX4 U377 ( .IN(n707), .OUT(n710) );
  INVX4 U378 ( .IN(Final_Exponent_reg[3]), .OUT(n407) );
  NANDX2 U379 ( .IN1(n946), .IN2(n912), .OUT(n235) );
  BUF4X U380 ( .IN(n1081), .OUT(Dataout_valid) );
  NANDX2 U381 ( .IN1(n235), .IN2(n236), .OUT(n230) );
  INVX4 U382 ( .IN(n1035), .OUT(n432) );
  BUF4X U383 ( .IN(n1059), .OUT(n402) );
  NAND2X1 U384 ( .IN1(C1_DATA9_0), .IN2(n818), .OUT(n507) );
  NAND2X1 U385 ( .IN1(n288), .IN2(n676), .OUT(n677) );
  NANDX2 U386 ( .IN1(n927), .IN2(n926), .OUT(n375) );
  NANDX2 U387 ( .IN1(n914), .IN2(n228), .OUT(n227) );
  NANDX2 U388 ( .IN1(n659), .IN2(n722), .OUT(n293) );
  NANDX2 U389 ( .IN1(n709), .IN2(n708), .OUT(n725) );
  INVX4 U390 ( .IN(n970), .OUT(n1009) );
  NANDX2 U391 ( .IN1(n409), .IN2(n946), .OUT(n301) );
  NAND2X1 U392 ( .IN1(Multi_dataout[10]), .IN2(n960), .OUT(n228) );
  NANDX2 U393 ( .IN1(n409), .IN2(n518), .OUT(n956) );
  INVX1 U394 ( .IN(n570), .OUT(n571) );
  NANDX2 U395 ( .IN1(n409), .IN2(n352), .OUT(n351) );
  NAND2X1 U396 ( .IN1(n299), .IN2(n960), .OUT(n290) );
  INVX1 U397 ( .IN(n287), .OUT(n286) );
  NANDX2 U398 ( .IN1(n880), .IN2(n879), .OUT(n959) );
  NANDX2 U399 ( .IN1(n457), .IN2(n549), .OUT(n1024) );
  INVX4 U400 ( .IN(n759), .OUT(n760) );
  NANDX2 U401 ( .IN1(n401), .IN2(n965), .OUT(n759) );
  NAND2X1 U402 ( .IN1(n599), .IN2(n781), .OUT(n600) );
  NAND2X1 U403 ( .IN1(DP_OP_343_164_2358_n38), .IN2(DP_OP_343_164_2358_n27), 
        .OUT(DP_OP_343_164_2358_n25) );
  NANDX2 U404 ( .IN1(n355), .IN2(n351), .OUT(n96) );
  NAND2X1 U405 ( .IN1(n782), .IN2(n781), .OUT(n784) );
  INVX1 U406 ( .IN(n768), .OUT(n769) );
  INVX1 U407 ( .IN(n766), .OUT(n767) );
  NAND2X1 U408 ( .IN1(Datain1[13]), .IN2(n411), .OUT(n384) );
  NANDX2 U409 ( .IN1(n867), .IN2(n866), .OUT(n868) );
  NAND2X1 U410 ( .IN1(n286), .IN2(n334), .OUT(n864) );
  NAND2X1 U411 ( .IN1(StateMC_0_), .IN2(n186), .OUT(n1036) );
  NANDX2 U412 ( .IN1(n409), .IN2(n945), .OUT(n740) );
  INVX4 U413 ( .IN(n541), .OUT(n660) );
  NANDX2 U414 ( .IN1(n494), .IN2(n659), .OUT(n721) );
  NAND2X1 U415 ( .IN1(n404), .IN2(Dataout_valid), .OUT(n1002) );
  NANDX2 U416 ( .IN1(n752), .IN2(n751), .OUT(n965) );
  INVX1 U417 ( .IN(DP_OP_345_166_2358_n35), .OUT(DP_OP_345_166_2358_n19) );
  INVX1 U418 ( .IN(DP_OP_348_169_2358_n31), .OUT(DP_OP_348_169_2358_n19) );
  NAND2X1 U419 ( .IN1(C1_DATA13_7), .IN2(n835), .OUT(n612) );
  INVX4 U420 ( .IN(n333), .OUT(n332) );
  NANDX2 U421 ( .IN1(n945), .IN2(n886), .OUT(n354) );
  INVX4 U422 ( .IN(n964), .OUT(n341) );
  NANDX2 U423 ( .IN1(n409), .IN2(n552), .OUT(n360) );
  NANDX2 U424 ( .IN1(n409), .IN2(n545), .OUT(n569) );
  INVX1 U425 ( .IN(DP_OP_340_161_2358_n11), .OUT(DP_OP_340_161_2358_n29) );
  INVX1 U426 ( .IN(DP_OP_340_161_2358_n15), .OUT(DP_OP_340_161_2358_n30) );
  INVX4 U427 ( .IN(n658), .OUT(n818) );
  INVX1 U428 ( .IN(DP_OP_341_162_2358_n15), .OUT(DP_OP_341_162_2358_n34) );
  INVX1 U429 ( .IN(DP_OP_341_162_2358_n23), .OUT(DP_OP_341_162_2358_n36) );
  INVX1 U430 ( .IN(DP_OP_339_160_2358_n23), .OUT(DP_OP_339_160_2358_n36) );
  INVX1 U431 ( .IN(DP_OP_339_160_2358_n27), .OUT(DP_OP_339_160_2358_n37) );
  NAND2X1 U432 ( .IN1(C1_DATA13_8), .IN2(n835), .OUT(n836) );
  INVX4 U433 ( .IN(n378), .OUT(n377) );
  NANDX2 U434 ( .IN1(Datain2[8]), .IN2(Datain1[8]), .OUT(n389) );
  NANDX2 U435 ( .IN1(n1012), .IN2(n735), .OUT(n543) );
  INVX4 U436 ( .IN(n283), .OUT(n282) );
  NAND2X1 U437 ( .IN1(Multi_dataout[6]), .IN2(n163), .OUT(n244) );
  NANDX2 U438 ( .IN1(n942), .IN2(n925), .OUT(n211) );
  NANDX2 U439 ( .IN1(n942), .IN2(n913), .OUT(n236) );
  INVX4 U440 ( .IN(n873), .OUT(n259) );
  NANDX2 U441 ( .IN1(n872), .IN2(n950), .OUT(n873) );
  INVX4 U442 ( .IN(n868), .OUT(n871) );
  INVX4 U443 ( .IN(n551), .OUT(n1013) );
  NANDX2 U444 ( .IN1(n531), .IN2(n738), .OUT(n532) );
  INVX4 U445 ( .IN(n413), .OUT(n420) );
  INVX4 U446 ( .IN(Datain2[13]), .OUT(n411) );
  INVX4 U447 ( .IN(Datain2[8]), .OUT(n412) );
  INVX4 U448 ( .IN(n424), .OUT(n430) );
  NAND2X1 U449 ( .IN1(n234), .IN2(n233), .OUT(n232) );
  INVX4 U450 ( .IN(n372), .OUT(n679) );
  NANDX2 U451 ( .IN1(n720), .IN2(n293), .OUT(n372) );
  INVX4 U452 ( .IN(n266), .OUT(n265) );
  NANDX2 U453 ( .IN1(n732), .IN2(n673), .OUT(n266) );
  INVX4 U454 ( .IN(n329), .OUT(n328) );
  NANDX2 U455 ( .IN1(n161), .IN2(n276), .OUT(n275) );
  INVX4 U456 ( .IN(n309), .OUT(n308) );
  INVX4 U457 ( .IN(n224), .OUT(n223) );
  NANDX2 U458 ( .IN1(n732), .IN2(n717), .OUT(n224) );
  NANDX2 U459 ( .IN1(n499), .IN2(n661), .OUT(n500) );
  NAND2X1 U460 ( .IN1(n466), .IN2(n307), .OUT(n346) );
  INVX4 U461 ( .IN(n668), .OUT(n481) );
  INVX4 U462 ( .IN(n1040), .OUT(n1012) );
  INVX4 U463 ( .IN(n862), .OUT(n731) );
  NANDX2 U464 ( .IN1(n728), .IN2(n268), .OUT(n862) );
  INVX4 U465 ( .IN(Multi_dataout[10]), .OUT(n209) );
  INVX4 U466 ( .IN(n368), .OUT(n367) );
  NANDX2 U467 ( .IN1(n409), .IN2(n1034), .OUT(n970) );
  NANDX2 U468 ( .IN1(n1040), .IN2(n409), .OUT(n1062) );
  NANDX2 U469 ( .IN1(n789), .IN2(N368), .OUT(n453) );
  NANDX2 U470 ( .IN1(n966), .IN2(n760), .OUT(n792) );
  INVX4 U471 ( .IN(n512), .OUT(n513) );
  NANDX2 U472 ( .IN1(n511), .IN2(n510), .OUT(n512) );
  INVX4 U473 ( .IN(n626), .OUT(n627) );
  NANDX2 U474 ( .IN1(n625), .IN2(n624), .OUT(n626) );
  INVX4 U475 ( .IN(n644), .OUT(n645) );
  NANDX2 U476 ( .IN1(n643), .IN2(n642), .OUT(n644) );
  INVX4 U477 ( .IN(n560), .OUT(n561) );
  NANDX2 U478 ( .IN1(n559), .IN2(n558), .OUT(n560) );
  NANDX2 U479 ( .IN1(n436), .IN2(n1043), .OUT(n1030) );
  NANDX2 U480 ( .IN1(n332), .IN2(n331), .OUT(n698) );
  NANDX2 U481 ( .IN1(n822), .IN2(C1_DATA2_7), .OUT(n364) );
  NANDX2 U482 ( .IN1(n354), .IN2(n353), .OUT(n352) );
  INVX4 U483 ( .IN(n340), .OUT(n339) );
  NANDX2 U484 ( .IN1(n341), .IN2(n362), .OUT(n340) );
  NANDX2 U485 ( .IN1(n888), .IN2(n889), .OUT(n963) );
  NANDX2 U486 ( .IN1(n748), .IN2(n306), .OUT(n886) );
  NANDX2 U487 ( .IN1(n357), .IN2(n788), .OUT(n356) );
  INVX4 U488 ( .IN(n358), .OUT(n357) );
  NANDX2 U489 ( .IN1(n850), .IN2(n841), .OUT(n358) );
  INVX4 U490 ( .IN(n360), .OUT(n359) );
  NANDX2 U491 ( .IN1(n184), .IN2(DP_OP_339_160_2358_n33), .OUT(n336) );
  INVX4 U492 ( .IN(n910), .OUT(n894) );
  NANDX2 U493 ( .IN1(n377), .IN2(n376), .OUT(n89) );
  NANDX2 U494 ( .IN1(n409), .IN2(n872), .OUT(n653) );
  INVX4 U495 ( .IN(DP_OP_347_168_2358_n38), .OUT(DP_OP_347_168_2358_n31) );
  NANDX2 U496 ( .IN1(n175), .IN2(DP_OP_345_166_2358_n23), .OUT(
        DP_OP_345_166_2358_n35) );
  INVX4 U497 ( .IN(DP_OP_345_166_2358_n36), .OUT(DP_OP_345_166_2358_n23) );
  NANDX2 U498 ( .IN1(n165), .IN2(n468), .OUT(DP_OP_345_166_2358_n36) );
  INVX4 U499 ( .IN(n714), .OUT(n821) );
  NANDX2 U500 ( .IN1(n175), .IN2(DP_OP_343_164_2358_n23), .OUT(n398) );
  NANDX2 U501 ( .IN1(n175), .IN2(DP_OP_340_161_2358_n23), .OUT(
        DP_OP_340_161_2358_n31) );
  INVX4 U502 ( .IN(DP_OP_340_161_2358_n32), .OUT(DP_OP_340_161_2358_n23) );
  NANDX2 U503 ( .IN1(n165), .IN2(DP_OP_340_161_2358_n27), .OUT(
        DP_OP_340_161_2358_n32) );
  NANDX2 U504 ( .IN1(n185), .IN2(DP_OP_349_170_2358_n19), .OUT(
        DP_OP_349_170_2358_n34) );
  INVX4 U505 ( .IN(DP_OP_349_170_2358_n35), .OUT(DP_OP_349_170_2358_n19) );
  NANDX2 U506 ( .IN1(n175), .IN2(DP_OP_349_170_2358_n23), .OUT(
        DP_OP_349_170_2358_n35) );
  NANDX2 U507 ( .IN1(n817), .IN2(C1_DATA4_8), .OUT(n318) );
  NANDX2 U508 ( .IN1(n175), .IN2(DP_OP_342_163_2358_n23), .OUT(n382) );
  INVX4 U509 ( .IN(DP_OP_342_163_2358_n28), .OUT(DP_OP_342_163_2358_n23) );
  INVX4 U510 ( .IN(n713), .OUT(n817) );
  INVX4 U511 ( .IN(n670), .OUT(n820) );
  NANDX2 U512 ( .IN1(n185), .IN2(DP_OP_351_172_2358_n19), .OUT(
        DP_OP_351_172_2358_n34) );
  INVX4 U513 ( .IN(DP_OP_351_172_2358_n35), .OUT(DP_OP_351_172_2358_n19) );
  NANDX2 U514 ( .IN1(n175), .IN2(DP_OP_351_172_2358_n23), .OUT(
        DP_OP_351_172_2358_n35) );
  INVX4 U515 ( .IN(n729), .OUT(n833) );
  INVX4 U516 ( .IN(n733), .OUT(n834) );
  NANDX2 U517 ( .IN1(n175), .IN2(DP_OP_348_169_2358_n23), .OUT(
        DP_OP_348_169_2358_n31) );
  INVX4 U518 ( .IN(n268), .OUT(n831) );
  NANDX2 U519 ( .IN1(n184), .IN2(DP_OP_344_165_2358_n15), .OUT(
        DP_OP_344_165_2358_n29) );
  INVX4 U520 ( .IN(DP_OP_344_165_2358_n30), .OUT(DP_OP_344_165_2358_n15) );
  NANDX2 U521 ( .IN1(n185), .IN2(DP_OP_344_165_2358_n19), .OUT(
        DP_OP_344_165_2358_n30) );
  INVX4 U522 ( .IN(n712), .OUT(n832) );
  INVX4 U523 ( .IN(n788), .OUT(N368) );
  INVX4 U524 ( .IN(n431), .OUT(RSOP_340_C1_Z_0) );
  NANDX2 U525 ( .IN1(n968), .IN2(n971), .OUT(n431) );
  INVX4 U526 ( .IN(n389), .OUT(DP_OP_269_159_6943_n102) );
  INVX4 U527 ( .IN(n388), .OUT(DP_OP_269_159_6943_n100) );
  NANDX2 U528 ( .IN1(n383), .IN2(n384), .OUT(DP_OP_269_159_6943_n93) );
  INVX4 U529 ( .IN(n385), .OUT(DP_OP_269_159_6943_n94) );
  INVX4 U530 ( .IN(n387), .OUT(DP_OP_269_159_6943_n98) );
  INVX4 U531 ( .IN(n386), .OUT(DP_OP_269_159_6943_n96) );
  NANDX2 U532 ( .IN1(n409), .IN2(n789), .OUT(n619) );
  INVX4 U533 ( .IN(n845), .OUT(n789) );
  NANDX2 U534 ( .IN1(n751), .IN2(n545), .OUT(n841) );
  NANDX2 U535 ( .IN1(n452), .IN2(n805), .OUT(n545) );
  NANDX2 U536 ( .IN1(n401), .IN2(n752), .OUT(n452) );
  INVX4 U537 ( .IN(n849), .OUT(n751) );
  NANDX2 U538 ( .IN1(n880), .IN2(n239), .OUT(n816) );
  INVX4 U539 ( .IN(n543), .OUT(n242) );
  INVX4 U540 ( .IN(n954), .OUT(n752) );
  INVX4 U541 ( .IN(n953), .OUT(n451) );
  NANDX2 U542 ( .IN1(n291), .IN2(n290), .OUT(n289) );
  INVX4 U543 ( .IN(n292), .OUT(n291) );
  NANDX2 U544 ( .IN1(n282), .IN2(n279), .OUT(n292) );
  NANDX2 U545 ( .IN1(n210), .IN2(n943), .OUT(n944) );
  NANDX2 U546 ( .IN1(n305), .IN2(n304), .OUT(n941) );
  NANDX2 U547 ( .IN1(n213), .IN2(n212), .OUT(n925) );
  NANDX2 U548 ( .IN1(n218), .IN2(n217), .OUT(n294) );
  NANDX2 U549 ( .IN1(n258), .IN2(n255), .OUT(n913) );
  INVX4 U550 ( .IN(n277), .OUT(n942) );
  NANDX2 U551 ( .IN1(n874), .IN2(n259), .OUT(n277) );
  NANDX2 U552 ( .IN1(n871), .IN2(n870), .OUT(n950) );
  INVX4 U553 ( .IN(n930), .OUT(n872) );
  NANDX2 U554 ( .IN1(n248), .IN2(n247), .OUT(n912) );
  INVX4 U555 ( .IN(n940), .OUT(n271) );
  NANDX2 U556 ( .IN1(n237), .IN2(n744), .OUT(n940) );
  INVX4 U557 ( .IN(n958), .OUT(n922) );
  INVX4 U558 ( .IN(n603), .OUT(n782) );
  INVX4 U559 ( .IN(n649), .OUT(n599) );
  NANDX2 U560 ( .IN1(DP_OP_349_170_2358_n55), .IN2(n650), .OUT(n649) );
  INVX4 U561 ( .IN(n468), .OUT(n650) );
  INVX4 U562 ( .IN(n401), .OUT(n921) );
  INVX4 U563 ( .IN(n933), .OUT(n924) );
  INVX4 U564 ( .IN(n520), .OUT(n957) );
  NANDX2 U565 ( .IN1(n755), .IN2(n519), .OUT(n938) );
  NANDX2 U566 ( .IN1(n528), .IN2(n1013), .OUT(n519) );
  NANDX2 U567 ( .IN1(n446), .IN2(n1013), .OUT(n755) );
  INVX4 U568 ( .IN(n956), .OUT(n916) );
  INVX4 U569 ( .IN(n936), .OUT(n518) );
  NANDX2 U570 ( .IN1(n528), .IN2(n517), .OUT(n936) );
  INVX4 U571 ( .IN(n532), .OUT(n844) );
  INVX4 U572 ( .IN(n445), .OUT(n987) );
  INVX4 U573 ( .IN(n457), .OUT(n528) );
  NANDX2 U574 ( .IN1(n1017), .IN2(n435), .OUT(n457) );
  INVX4 U575 ( .IN(n438), .OUT(n988) );
  NANDX2 U576 ( .IN1(n801), .IN2(n757), .OUT(n845) );
  NANDX2 U577 ( .IN1(n420), .IN2(n419), .OUT(n968) );
  NANDX2 U578 ( .IN1(n430), .IN2(n429), .OUT(n971) );
  INVX4 U579 ( .IN(Datain1[11]), .OUT(n426) );
  INVX4 U580 ( .IN(Datain1[10]), .OUT(n427) );
  INVX4 U581 ( .IN(Datain1[13]), .OUT(n422) );
  INVX4 U582 ( .IN(Datain1[8]), .OUT(n423) );
  NANDX2 U583 ( .IN1(n249), .IN2(n237), .OUT(n251) );
  INVX4 U584 ( .IN(n243), .OUT(n237) );
  NANDX2 U585 ( .IN1(n249), .IN2(n164), .OUT(n219) );
  NANDX2 U586 ( .IN1(n744), .IN2(n164), .OUT(n295) );
  NANDX2 U587 ( .IN1(n265), .IN2(n260), .OUT(n243) );
  NANDX2 U588 ( .IN1(n675), .IN2(n674), .OUT(n678) );
  NANDX2 U589 ( .IN1(n315), .IN2(n317), .OUT(n672) );
  INVX4 U590 ( .IN(n316), .OUT(n315) );
  NANDX2 U591 ( .IN1(n670), .IN2(n714), .OUT(n316) );
  INVX4 U592 ( .IN(n249), .OUT(n744) );
  NANDX2 U593 ( .IN1(n669), .IN2(n267), .OUT(n249) );
  NANDX2 U594 ( .IN1(n701), .IN2(n495), .OUT(n664) );
  INVX4 U595 ( .IN(n700), .OUT(n495) );
  NANDX2 U596 ( .IN1(n348), .IN2(n939), .OUT(n700) );
  INVX4 U597 ( .IN(n349), .OUT(n348) );
  NANDX2 U598 ( .IN1(n269), .IN2(n661), .OUT(n701) );
  INVX4 U599 ( .IN(n270), .OUT(n269) );
  NANDX2 U600 ( .IN1(n663), .IN2(n662), .OUT(n675) );
  INVX4 U601 ( .IN(n275), .OUT(n274) );
  NANDX2 U602 ( .IN1(n498), .IN2(n497), .OUT(n658) );
  INVX4 U603 ( .IN(n505), .OUT(n663) );
  NANDX2 U604 ( .IN1(n739), .IN2(n874), .OUT(n911) );
  NANDX2 U605 ( .IN1(n223), .IN2(n221), .OUT(n947) );
  NANDX2 U606 ( .IN1(n394), .IN2(n222), .OUT(n221) );
  INVX4 U607 ( .IN(n537), .OUT(n718) );
  NANDX2 U608 ( .IN1(n706), .IN2(n484), .OUT(n712) );
  NANDX2 U609 ( .IN1(n403), .IN2(n483), .OUT(n705) );
  NANDX2 U610 ( .IN1(n482), .IN2(n661), .OUT(n706) );
  NANDX2 U611 ( .IN1(n504), .IN2(n702), .OUT(n714) );
  INVX4 U612 ( .IN(n666), .OUT(n504) );
  NANDX2 U613 ( .IN1(n500), .IN2(n505), .OUT(n666) );
  NANDX2 U614 ( .IN1(n406), .IN2(n661), .OUT(n505) );
  NANDX2 U615 ( .IN1(n475), .IN2(n474), .OUT(n711) );
  INVX4 U616 ( .IN(n676), .OUT(n474) );
  NANDX2 U617 ( .IN1(n473), .IN2(n483), .OUT(n676) );
  INVX4 U618 ( .IN(n493), .OUT(n661) );
  NANDX2 U619 ( .IN1(n394), .IN2(DP_OP_341_162_2358_n38), .OUT(n468) );
  NANDX2 U620 ( .IN1(n733), .IN2(n732), .OUT(n869) );
  NANDX2 U621 ( .IN1(n369), .IN2(n865), .OUT(n732) );
  INVX4 U622 ( .IN(n724), .OUT(n865) );
  NANDX2 U623 ( .IN1(n347), .IN2(n220), .OUT(n724) );
  INVX4 U624 ( .IN(n476), .OUT(n499) );
  NANDX2 U625 ( .IN1(n491), .IN2(n722), .OUT(n733) );
  INVX4 U626 ( .IN(n490), .OUT(n722) );
  NANDX2 U627 ( .IN1(n326), .IN2(n347), .OUT(n490) );
  INVX4 U628 ( .IN(n327), .OUT(n326) );
  NANDX2 U629 ( .IN1(n307), .IN2(Multi_dataout[1]), .OUT(n327) );
  INVX4 U630 ( .IN(Multi_dataout[2]), .OUT(n307) );
  INVX4 U631 ( .IN(n659), .OUT(n491) );
  NANDX2 U632 ( .IN1(n731), .IN2(n730), .OUT(n734) );
  NANDX2 U633 ( .IN1(n481), .IN2(n667), .OUT(n317) );
  INVX4 U634 ( .IN(n288), .OUT(n667) );
  NANDX2 U635 ( .IN1(n480), .IN2(n492), .OUT(n288) );
  NANDX2 U636 ( .IN1(n803), .IN2(n458), .OUT(n930) );
  NANDX2 U637 ( .IN1(n1012), .IN2(Multi_ack), .OUT(n810) );
  INVX4 U638 ( .IN(n433), .OUT(n1014) );
  NAND2X1 U639 ( .IN1(n180), .IN2(n179), .OUT(n433) );
  NANDX2 U640 ( .IN1(n489), .IN2(n708), .OUT(n268) );
  INVX4 U641 ( .IN(n863), .OUT(n708) );
  NANDX2 U642 ( .IN1(n488), .IN2(n182), .OUT(n863) );
  INVX4 U643 ( .IN(n535), .OUT(n472) );
  INVX4 U644 ( .IN(n478), .OUT(n502) );
  NANDX2 U645 ( .IN1(n209), .IN2(n470), .OUT(n478) );
  NANDX2 U646 ( .IN1(n367), .IN2(n347), .OUT(n728) );
  NANDX2 U647 ( .IN1(n322), .IN2(n321), .OUT(n467) );
  NANDX2 U648 ( .IN1(n350), .IN2(n477), .OUT(n486) );
  INVX4 U649 ( .IN(n390), .OUT(n477) );
  INVX4 U650 ( .IN(n391), .OUT(n350) );
  INVX4 U651 ( .IN(Multi_dataout[11]), .OUT(n470) );
  INVX4 U652 ( .IN(n323), .OUT(n322) );
  NANDX2 U653 ( .IN1(n325), .IN2(n324), .OUT(n323) );
  NANDX2 U654 ( .IN1(n399), .IN2(n903), .OUT(n535) );
  INVX4 U655 ( .IN(Multi_dataout[8]), .OUT(n903) );
  INVX4 U656 ( .IN(Multi_dataout[9]), .OUT(n399) );
  INVX4 U657 ( .IN(n463), .OUT(n325) );
  NANDX2 U658 ( .IN1(n471), .IN2(n469), .OUT(n463) );
  INVX4 U659 ( .IN(Multi_dataout[6]), .OUT(n469) );
  INVX4 U660 ( .IN(Multi_dataout[12]), .OUT(n471) );
  NANDX2 U661 ( .IN1(n406), .IN2(n462), .OUT(n485) );
  INVX4 U662 ( .IN(Final_Exponent_reg[2]), .OUT(n406) );
  NANDX2 U663 ( .IN1(n407), .IN2(n462), .OUT(n493) );
  INVX4 U664 ( .IN(n461), .OUT(n462) );
  NANDX2 U665 ( .IN1(n392), .IN2(C1_DATA8_0), .OUT(DP_OP_345_166_2358_n31) );
  INVX4 U666 ( .IN(n392), .OUT(C1_DATA2_1) );
  INVX4 U667 ( .IN(RSTn_BAR), .OUT(n409) );
  INVX1 U668 ( .IN(Exc_Ack), .OUT(n809) );
  NAND2X1 U669 ( .IN1(Final_Mantissa_reg[0]), .IN2(Dataout_valid), .OUT(n994)
         );
  NAND2X1 U670 ( .IN1(Final_Mantissa_reg[1]), .IN2(Dataout_valid), .OUT(n995)
         );
  NAND2X1 U671 ( .IN1(Final_Mantissa_reg[2]), .IN2(Dataout_valid), .OUT(n996)
         );
  NAND2X1 U672 ( .IN1(Final_Mantissa_reg[3]), .IN2(Dataout_valid), .OUT(n997)
         );
  NAND2X1 U673 ( .IN1(DP_OP_349_170_2358_n56), .IN2(Dataout_valid), .OUT(n1005) );
  INVX1 U674 ( .IN(Dataout_valid), .OUT(n1031) );
  NAND2X1 U675 ( .IN1(n394), .IN2(Dataout_valid), .OUT(n1003) );
  NAND2X1 U676 ( .IN1(DP_OP_349_170_2358_n57), .IN2(Dataout_valid), .OUT(n1006) );
  NAND2X1 U677 ( .IN1(Final_Mantissa_reg[4]), .IN2(Dataout_valid), .OUT(n998)
         );
  NAND2X1 U678 ( .IN1(DP_OP_349_170_2358_n55), .IN2(Dataout_valid), .OUT(n1004) );
  NAND2X1 U679 ( .IN1(DP_OP_349_170_2358_n58), .IN2(Dataout_valid), .OUT(n1007) );
  NAND2X1 U680 ( .IN1(n181), .IN2(Dataout_valid), .OUT(n1008) );
  NAND2X1 U681 ( .IN1(Final_Mantissa_reg[6]), .IN2(Dataout_valid), .OUT(n1000)
         );
  INVX1 U682 ( .IN(n971), .OUT(n967) );
  INVX1 U683 ( .IN(n965), .OUT(n1025) );
  NAND2X1 U684 ( .IN1(n409), .IN2(n455), .OUT(n417) );
  NAND2X1 U685 ( .IN1(Exc_value[1]), .IN2(n791), .OUT(n448) );
  INVX1 U686 ( .IN(n765), .OUT(n405) );
  NAND2X1 U687 ( .IN1(n991), .IN2(n755), .OUT(n756) );
  NAND2X1 U688 ( .IN1(n200), .IN2(Dataout_valid), .OUT(n991) );
  INVX1 U689 ( .IN(n798), .OUT(n521) );
  NAND2X1 U690 ( .IN1(n993), .IN2(n850), .OUT(n790) );
  NAND2X1 U691 ( .IN1(n193), .IN2(Dataout_valid), .OUT(n993) );
  NAND2X1 U692 ( .IN1(Exc_Ack), .IN2(n1010), .OUT(n447) );
  NAND2X1 U693 ( .IN1(n1012), .IN2(n750), .OUT(n753) );
  INVX1 U694 ( .IN(DP_OP_348_169_2358_n23), .OUT(DP_OP_348_169_2358_n32) );
  NAND2X1 U695 ( .IN1(DP_OP_341_162_2358_n38), .IN2(n781), .OUT(n634) );
  INVX1 U696 ( .IN(n785), .OUT(n654) );
  NAND2X1 U697 ( .IN1(C1_DATA13_5), .IN2(n835), .OUT(n575) );
  INVX1 U698 ( .IN(DP_OP_351_172_2358_n34), .OUT(DP_OP_351_172_2358_n15) );
  INVX1 U699 ( .IN(DP_OP_349_170_2358_n34), .OUT(DP_OP_349_170_2358_n15) );
  INVX1 U700 ( .IN(n808), .OUT(n548) );
  INVX1 U701 ( .IN(n526), .OUT(n434) );
  INVX1 U702 ( .IN(n757), .OUT(n758) );
  INVX1 U703 ( .IN(n606), .OUT(n607) );
  NAND2X1 U704 ( .IN1(n409), .IN2(Multi_dataout[13]), .OUT(n296) );
  NAND2X1 U705 ( .IN1(n947), .IN2(n948), .OUT(n362) );
  NAND2X1 U706 ( .IN1(n343), .IN2(n748), .OUT(n342) );
  INVX1 U707 ( .IN(n887), .OUT(n343) );
  NAND2X1 U708 ( .IN1(n874), .IN2(n306), .OUT(n361) );
  NAND2X1 U709 ( .IN1(n962), .IN2(n961), .OUT(n381) );
  NAND2X1 U710 ( .IN1(Datain1[2]), .IN2(n916), .OUT(n891) );
  NAND2X1 U711 ( .IN1(n409), .IN2(n942), .OUT(n900) );
  INVX1 U712 ( .IN(n238), .OUT(n783) );
  NAND2X1 U713 ( .IN1(C1_DATA13_6), .IN2(n835), .OUT(n773) );
  INVX1 U714 ( .IN(Datain1[0]), .OUT(n851) );
  INVX1 U715 ( .IN(n403), .OUT(n854) );
  INVX1 U716 ( .IN(n959), .OUT(n882) );
  NAND2X1 U717 ( .IN1(n393), .IN2(n190), .OUT(DP_OP_347_168_2358_n38) );
  NAND2X1 U718 ( .IN1(n166), .IN2(n407), .OUT(DP_OP_342_163_2358_n28) );
  NAND2X1 U719 ( .IN1(Datain2[9]), .IN2(Datain1[9]), .OUT(n388) );
  NAND2X1 U720 ( .IN1(Datain2[13]), .IN2(n422), .OUT(n383) );
  NAND2X1 U721 ( .IN1(Datain2[12]), .IN2(Datain1[12]), .OUT(n385) );
  NAND2X1 U722 ( .IN1(Datain2[10]), .IN2(Datain1[10]), .OUT(n387) );
  NAND2X1 U723 ( .IN1(Datain2[11]), .IN2(Datain1[11]), .OUT(n386) );
  INVX1 U724 ( .IN(n841), .OUT(n380) );
  INVX1 U725 ( .IN(n816), .OUT(n843) );
  NAND2X1 U726 ( .IN1(n409), .IN2(Multi_dataout[12]), .OUT(n300) );
  NAND2X1 U727 ( .IN1(n932), .IN2(n947), .OUT(n284) );
  INVX1 U728 ( .IN(Datain1[5]), .OUT(n937) );
  NAND2X1 U729 ( .IN1(Multi_dataout[0]), .IN2(n170), .OUT(n258) );
  INVX1 U730 ( .IN(n869), .OUT(n870) );
  NAND2X1 U731 ( .IN1(n346), .IN2(n347), .OUT(n334) );
  NAND2X1 U732 ( .IN1(n288), .IN2(n863), .OUT(n287) );
  INVX1 U733 ( .IN(Multi_dataout[15]), .OUT(n735) );
  NAND2X1 U734 ( .IN1(n849), .IN2(n848), .OUT(n958) );
  NAND2X1 U735 ( .IN1(Final_Mantissa_reg[2]), .IN2(n890), .OUT(n907) );
  NAND2X1 U736 ( .IN1(Exc_Ack), .IN2(n988), .OUT(n812) );
  NAND2X1 U737 ( .IN1(n409), .IN2(n878), .OUT(n879) );
  NAND2X1 U738 ( .IN1(n845), .IN2(n844), .OUT(n878) );
  NAND2X1 U739 ( .IN1(Exc_Ack), .IN2(n1024), .OUT(n529) );
  NAND2X1 U740 ( .IN1(Exc_Ack), .IN2(n528), .OUT(n530) );
  INVX1 U741 ( .IN(Exc_value[0]), .OUT(n435) );
  INVX1 U742 ( .IN(Exc_value[2]), .OUT(n1016) );
  INVX1 U743 ( .IN(Datain2[14]), .OUT(n415) );
  INVX1 U744 ( .IN(Datain2[7]), .OUT(n416) );
  NAND2X1 U745 ( .IN1(n192), .IN2(n1014), .OUT(n526) );
  NAND2X1 U746 ( .IN1(n409), .IN2(n401), .OUT(n952) );
  BUF4X U747 ( .IN(n1011), .OUT(n401) );
  NAND2X1 U748 ( .IN1(C1_DATA2_1), .IN2(n664), .OUT(n329) );
  NAND2X1 U749 ( .IN1(n406), .IN2(C1_DATA2_1), .OUT(n270) );
  INVX1 U750 ( .IN(n533), .OUT(n534) );
  NAND2X1 U751 ( .IN1(n661), .IN2(n391), .OUT(n309) );
  INVX1 U752 ( .IN(n721), .OUT(n723) );
  NAND2X1 U753 ( .IN1(n394), .IN2(n392), .OUT(n482) );
  NAND2X1 U754 ( .IN1(n733), .IN2(n711), .OUT(n716) );
  INVX4 U755 ( .IN(n166), .OUT(n394) );
  INVX1 U756 ( .IN(Multi_dataout[3]), .OUT(n487) );
  BUF4X U757 ( .IN(Multi_dataout[4]), .OUT(n390) );
  NAND2X1 U758 ( .IN1(Multi_dataout[2]), .IN2(n721), .OUT(n368) );
  INVX4 U759 ( .IN(C1_DATA2_1), .OUT(n404) );
  BUF4X U760 ( .IN(Final_Exponent_reg[1]), .OUT(n392) );
  INVX4 U761 ( .IN(n183), .OUT(DP_OP_349_170_2358_n56) );
  INVX4 U762 ( .IN(n185), .OUT(DP_OP_349_170_2358_n57) );
  INVX1 U763 ( .IN(Multi_dataout[1]), .OUT(n466) );
  INVX4 U764 ( .IN(n184), .OUT(DP_OP_349_170_2358_n58) );
  INVX1 U765 ( .IN(Multi_dataout[0]), .OUT(n931) );
  INVX4 U766 ( .IN(n189), .OUT(n408) );
  AOI22 U767 ( .IN1(n168), .IN2(Multi_dataout[2]), .IN3(n271), .IN4(
        Multi_dataout[3]), .OUT(n212) );
  AOI22 U768 ( .IN1(n278), .IN2(Multi_dataout[0]), .IN3(Multi_dataout[1]), 
        .IN4(n170), .OUT(n213) );
  AOI22 U769 ( .IN1(n168), .IN2(Multi_dataout[6]), .IN3(n271), .IN4(n403), 
        .OUT(n217) );
  AOI22 U770 ( .IN1(n278), .IN2(n390), .IN3(n391), .IN4(n170), .OUT(n218) );
  AOI22 U771 ( .IN1(n278), .IN2(Multi_dataout[3]), .IN3(n168), .IN4(n391), 
        .OUT(n248) );
  NOR2X1 U772 ( .IN1(n931), .IN2(n346), .OUT(n220) );
  INVX4 U773 ( .IN(n467), .OUT(n347) );
  NOR2X1 U774 ( .IN1(n369), .IN2(n724), .OUT(n370) );
  NAND3X1 U775 ( .IN1(n726), .IN2(n724), .IN3(n225), .OUT(n222) );
  INVX4 U776 ( .IN(n947), .OUT(n874) );
  NOR2X1 U777 ( .IN1(n226), .IN2(n727), .OUT(n225) );
  AOI22 U778 ( .IN1(n170), .IN2(n403), .IN3(Multi_dataout[8]), .IN4(n168), 
        .OUT(n889) );
  OAI21 U779 ( .IN1(n227), .IN2(n230), .IN3(n409), .OUT(n229) );
  AOI21 U780 ( .IN1(n171), .IN2(n232), .IN3(n906), .OUT(n231) );
  AOI22 U781 ( .IN1(n168), .IN2(n395), .IN3(n403), .IN4(n160), .OUT(n234) );
  NAND2X1 U782 ( .IN1(n237), .IN2(n297), .OUT(n257) );
  NOR2X1 U783 ( .IN1(n241), .IN2(n584), .OUT(n240) );
  MUX2X1 U784 ( .IN1(Multi_dataout[1]), .IN2(Multi_dataout[0]), .S(n164), 
        .OUT(n743) );
  INVX1 U785 ( .IN(Multi_dataout[13]), .OUT(n939) );
  NOR2X1 U786 ( .IN1(Multi_dataout[12]), .IN2(Multi_dataout[13]), .OUT(n501)
         );
  INVX4 U787 ( .IN(n746), .OUT(n946) );
  NAND3X1 U788 ( .IN1(n246), .IN2(n245), .IN3(n244), .OUT(n397) );
  AOI22 U789 ( .IN1(n278), .IN2(n391), .IN3(n403), .IN4(n168), .OUT(n245) );
  AOI22 U790 ( .IN1(n170), .IN2(n390), .IN3(Multi_dataout[6]), .IN4(n271), 
        .OUT(n247) );
  OAI21 U791 ( .IN1(n940), .IN2(n911), .IN3(n910), .OUT(n960) );
  NOR2X1 U792 ( .IN1(n307), .IN2(n249), .OUT(n297) );
  OAI21 U793 ( .IN1(n250), .IN2(n900), .IN3(n899), .OUT(n901) );
  AOI22 U794 ( .IN1(n168), .IN2(Multi_dataout[0]), .IN3(Multi_dataout[1]), 
        .IN4(n271), .OUT(n250) );
  OAI21 U795 ( .IN1(n399), .IN2(n251), .IN3(n915), .OUT(n920) );
  AOI22 U796 ( .IN1(Final_Mantissa_reg[0]), .IN2(n241), .IN3(n409), .IN4(n252), 
        .OUT(n363) );
  AOI21 U797 ( .IN1(n294), .IN2(n945), .IN3(n858), .OUT(n253) );
  OAI21 U798 ( .IN1(n295), .IN2(n466), .IN3(n257), .OUT(n256) );
  OAI21 U799 ( .IN1(n262), .IN2(n261), .IN3(C1_DATA8_0), .OUT(n260) );
  OAI21 U800 ( .IN1(n370), .IN2(n371), .IN3(n373), .OUT(n267) );
  AOI22 U801 ( .IN1(n278), .IN2(Multi_dataout[6]), .IN3(n395), .IN4(n271), 
        .OUT(n888) );
  NAND3X1 U802 ( .IN1(n293), .IN2(n274), .IN3(n272), .OUT(n371) );
  NOR2X1 U803 ( .IN1(n310), .IN2(n273), .OUT(n272) );
  NAND3X1 U804 ( .IN1(n950), .IN2(n281), .IN3(n280), .OUT(n279) );
  NOR2X1 U805 ( .IN1(RSTn_BAR), .IN2(n940), .OUT(n280) );
  AOI21 U806 ( .IN1(n397), .IN2(n172), .IN3(n289), .OUT(n302) );
  AOI22 U807 ( .IN1(n278), .IN2(Multi_dataout[1]), .IN3(Multi_dataout[3]), 
        .IN4(n168), .OUT(n305) );
  AOI22 U808 ( .IN1(n941), .IN2(n298), .IN3(n171), .IN4(n944), .OUT(n303) );
  AOI22 U809 ( .IN1(n271), .IN2(n390), .IN3(n170), .IN4(Multi_dataout[2]), 
        .OUT(n304) );
  AOI22 U810 ( .IN1(n160), .IN2(n395), .IN3(Multi_dataout[11]), .IN4(n168), 
        .OUT(n943) );
  AOI22 U811 ( .IN1(n278), .IN2(Multi_dataout[10]), .IN3(Multi_dataout[12]), 
        .IN4(n168), .OUT(n962) );
  AOI22 U812 ( .IN1(Multi_dataout[2]), .IN2(n278), .IN3(n390), .IN4(n168), 
        .OUT(n306) );
  AOI21 U813 ( .IN1(n702), .IN2(n666), .IN3(n665), .OUT(n311) );
  NOR2X1 U814 ( .IN1(n314), .IN2(n313), .OUT(n492) );
  NOR2X1 U815 ( .IN1(n158), .IN2(n314), .OUT(n483) );
  NAND2X1 U816 ( .IN1(Multi_dataout[3]), .IN2(n170), .OUT(n748) );
  OAI21 U817 ( .IN1(n320), .IN2(n319), .IN3(n318), .OUT(n819) );
  NOR2X1 U818 ( .IN1(n408), .IN2(DP_OP_341_162_2358_n3), .OUT(n319) );
  OAI21 U819 ( .IN1(n177), .IN2(DP_OP_341_162_2358_n3), .IN3(n818), .OUT(n320)
         );
  NOR2X1 U820 ( .IN1(n465), .IN2(n486), .OUT(n321) );
  NOR2X1 U821 ( .IN1(Multi_dataout[3]), .IN2(n535), .OUT(n324) );
  AOI22 U822 ( .IN1(n160), .IN2(Multi_dataout[8]), .IN3(Multi_dataout[10]), 
        .IN4(n168), .OUT(n915) );
  AOI21 U823 ( .IN1(n172), .IN2(n963), .IN3(n330), .OUT(n337) );
  OAI21 U824 ( .IN1(n615), .IN2(n616), .IN3(n951), .OUT(n331) );
  AOI22 U825 ( .IN1(n822), .IN2(C1_DATA2_6), .IN3(n336), .IN4(n335), .OUT(n768) );
  AOI21 U826 ( .IN1(DP_OP_339_160_2358_n15), .IN2(DP_OP_339_160_2358_n33), 
        .IN3(n670), .OUT(n335) );
  NAND3X1 U827 ( .IN1(n344), .IN2(n338), .IN3(n337), .OUT(n699) );
  OAI21 U828 ( .IN1(n361), .IN2(n342), .IN3(n339), .OUT(n338) );
  AOI21 U829 ( .IN1(n381), .IN2(n171), .IN3(n345), .OUT(n344) );
  INVX1 U830 ( .IN(n674), .OUT(n396) );
  NOR2X1 U831 ( .IN1(n350), .IN2(n940), .OUT(n887) );
  AOI21 U832 ( .IN1(n887), .IN2(n945), .IN3(n747), .OUT(n353) );
  NANDX2 U833 ( .IN1(n359), .IN2(n356), .OUT(n785) );
  NOR2X1 U834 ( .IN1(n887), .IN2(n886), .OUT(n949) );
  OAI21 U835 ( .IN1(n366), .IN2(n365), .IN3(n364), .OUT(n608) );
  NOR2X1 U836 ( .IN1(n181), .IN2(DP_OP_339_160_2358_n7), .OUT(n365) );
  OAI21 U837 ( .IN1(DP_OP_339_160_2358_n33), .IN2(DP_OP_339_160_2358_n7), 
        .IN3(n820), .OUT(n366) );
  OAI21 U838 ( .IN1(n375), .IN2(n374), .IN3(n409), .OUT(n928) );
  OAI21 U839 ( .IN1(n839), .IN2(n840), .IN3(n951), .OUT(n376) );
  OAI21 U840 ( .IN1(n189), .IN2(n843), .IN3(n379), .OUT(n378) );
  AOI22 U841 ( .IN1(n409), .IN2(n380), .IN3(n842), .IN4(N368), .OUT(n379) );
  NAND2X1 U842 ( .IN1(Final_Mantissa_reg[5]), .IN2(Dataout_valid), .OUT(n999)
         );
  INVX4 U843 ( .IN(n393), .OUT(C1_DATA8_0) );
  TIEHI U844 ( .OUT(n59) );
  NAND2X1 U845 ( .IN1(Multi_dataout[12]), .IN2(n939), .OUT(n538) );
  NAND2X1 U846 ( .IN1(n404), .IN2(DP_OP_345_166_2358_n31), .OUT(
        DP_OP_341_162_2358_n28) );
  NAND2X1 U847 ( .IN1(Final_Exponent_reg[0]), .IN2(DP_OP_345_166_2358_n31), 
        .OUT(DP_OP_341_162_2358_n29) );
  NAND2X1 U848 ( .IN1(C1_DATA2_1), .IN2(C1_DATA9_0), .OUT(n476) );
  NAND2X1 U849 ( .IN1(n535), .IN2(n534), .OUT(n536) );
  NAND2X1 U850 ( .IN1(C1_DATA8_0), .IN2(Dataout_valid), .OUT(n1001) );
  INVX1 U851 ( .IN(DP_OP_347_168_2358_n15), .OUT(DP_OP_347_168_2358_n34) );
  INVX1 U852 ( .IN(DP_OP_347_168_2358_n11), .OUT(DP_OP_347_168_2358_n33) );
  NAND2X1 U853 ( .IN1(n553), .IN2(n785), .OUT(n691) );
  NAND2X1 U854 ( .IN1(Multi_dataout[8]), .IN2(n399), .OUT(n503) );
  INVX1 U855 ( .IN(DP_OP_339_160_2358_n19), .OUT(DP_OP_339_160_2358_n35) );
  INVX1 U856 ( .IN(DP_OP_340_161_2358_n7), .OUT(DP_OP_340_161_2358_n28) );
  NAND2X1 U857 ( .IN1(Multi_dataout[11]), .IN2(n163), .OUT(n961) );
  INVX1 U858 ( .IN(DP_OP_343_164_2358_n23), .OUT(DP_OP_343_164_2358_n36) );
  INVX1 U859 ( .IN(n823), .OUT(n824) );
  INVX1 U860 ( .IN(DP_OP_343_164_2358_n7), .OUT(DP_OP_343_164_2358_n32) );
  INVX1 U861 ( .IN(DP_OP_341_162_2358_n11), .OUT(DP_OP_341_162_2358_n33) );
  INVX4 U862 ( .IN(n1061), .OUT(n1079) );
  NOR2X1 U863 ( .IN1(Datain2[9]), .IN2(Datain2[11]), .OUT(n410) );
  NAND3X1 U864 ( .IN1(n412), .IN2(n411), .IN3(n410), .OUT(n413) );
  NOR2X1 U865 ( .IN1(Datain2[10]), .IN2(Datain2[12]), .OUT(n414) );
  NAND3X1 U866 ( .IN1(n416), .IN2(n415), .IN3(n414), .OUT(n418) );
  NOR2X1 U867 ( .IN1(Datain1[12]), .IN2(Datain1[9]), .OUT(n421) );
  NAND3X1 U868 ( .IN1(n423), .IN2(n422), .IN3(n421), .OUT(n424) );
  NOR2X1 U869 ( .IN1(Datain1[14]), .IN2(Datain1[7]), .OUT(n425) );
  NAND3X1 U870 ( .IN1(n427), .IN2(n426), .IN3(n425), .OUT(n428) );
  NAND3X1 U871 ( .IN1(StateMC_0_), .IN2(n191), .IN3(n179), .OUT(n438) );
  OAI21 U872 ( .IN1(n528), .IN2(n809), .IN3(n988), .OUT(n436) );
  NOR2X1 U873 ( .IN1(n180), .IN2(n1036), .OUT(n1081) );
  NOR2X1 U874 ( .IN1(n180), .IN2(StateMC_0_), .OUT(n437) );
  NAND3X1 U875 ( .IN1(n445), .IN2(n438), .IN3(n990), .OUT(n439) );
  NOR2X1 U876 ( .IN1(Datain2[14]), .IN2(n971), .OUT(n443) );
  NAND3X1 U877 ( .IN1(Datain2[12]), .IN2(Datain2[7]), .IN3(n1023), .OUT(n442)
         );
  NOR2X1 U878 ( .IN1(Datain1[14]), .IN2(n968), .OUT(n441) );
  NAND3X1 U879 ( .IN1(Datain1[12]), .IN2(Datain1[7]), .IN3(n1020), .OUT(n440)
         );
  AOI22 U880 ( .IN1(n443), .IN2(n442), .IN3(n441), .IN4(n440), .OUT(n757) );
  NAND3X1 U881 ( .IN1(n1033), .IN2(n754), .IN3(n845), .OUT(n450) );
  NOR2X1 U882 ( .IN1(n206), .IN2(n205), .OUT(n444) );
  NAND3X1 U883 ( .IN1(Exc_value[0]), .IN2(Exc_value[1]), .IN3(n444), .OUT(n456) );
  NOR2X1 U884 ( .IN1(n550), .IN2(n456), .OUT(n446) );
  NAND3X1 U885 ( .IN1(n812), .IN2(n447), .IN3(n519), .OUT(n791) );
  NAND3X1 U886 ( .IN1(n755), .IN2(n992), .IN3(n448), .OUT(n449) );
  AOI21 U887 ( .IN1(n202), .IN2(n450), .IN3(n449), .OUT(n454) );
  MUX2X1 U888 ( .IN1(n408), .IN2(n189), .S(n605), .OUT(n849) );
  NOR2X1 U889 ( .IN1(n191), .IN2(n1036), .OUT(n1011) );
  INVX4 U890 ( .IN(n810), .OUT(n803) );
  NAND3X1 U891 ( .IN1(n454), .IN2(n841), .IN3(n453), .OUT(n455) );
  NOR2X1 U892 ( .IN1(Multi_dataout[15]), .IN2(Multi_dataout[14]), .OUT(n458)
         );
  NOR2X1 U893 ( .IN1(Final_Exponent_reg[4]), .IN2(Final_Exponent_reg[5]), 
        .OUT(n460) );
  NOR2X1 U894 ( .IN1(Final_Exponent_reg[6]), .IN2(Final_Exponent_reg[7]), 
        .OUT(n459) );
  NAND3X1 U895 ( .IN1(n189), .IN2(n460), .IN3(n459), .OUT(n461) );
  NOR2X1 U896 ( .IN1(Multi_dataout[10]), .IN2(n403), .OUT(n464) );
  NAND3X1 U897 ( .IN1(n470), .IN2(n939), .IN3(n464), .OUT(n465) );
  NOR2X1 U898 ( .IN1(n403), .IN2(n469), .OUT(n473) );
  OAI21 U899 ( .IN1(n476), .IN2(n485), .IN3(n493), .OUT(n668) );
  NOR2X1 U900 ( .IN1(n391), .IN2(n477), .OUT(n480) );
  NOR2X1 U901 ( .IN1(n403), .IN2(Multi_dataout[6]), .OUT(n479) );
  AOI22 U902 ( .IN1(n827), .IN2(C1_DATA9_0), .IN3(n826), .IN4(C1_DATA9_0), 
        .OUT(n515) );
  OAI21 U903 ( .IN1(n404), .IN2(n485), .IN3(n493), .OUT(n709) );
  NOR2X1 U904 ( .IN1(n487), .IN2(n486), .OUT(n488) );
  AOI22 U905 ( .IN1(n832), .IN2(C1_DATA8_0), .IN3(n831), .IN4(C1_DATA8_0), 
        .OUT(n514) );
  AOI22 U906 ( .IN1(n834), .IN2(Final_Exponent_reg[0]), .IN3(C1_DATA8_0), 
        .IN4(n833), .OUT(n511) );
  AOI22 U907 ( .IN1(n820), .IN2(C1_DATA9_0), .IN3(C1_DATA8_0), .IN4(n822), 
        .OUT(n508) );
  NOR2X1 U908 ( .IN1(n503), .IN2(n533), .OUT(n702) );
  NOR2X1 U909 ( .IN1(n399), .IN2(n533), .OUT(n662) );
  AOI22 U910 ( .IN1(n821), .IN2(C1_DATA9_0), .IN3(n817), .IN4(C1_DATA8_0), 
        .OUT(n506) );
  NAND3X1 U911 ( .IN1(n508), .IN2(n507), .IN3(n506), .OUT(n509) );
  AOI21 U912 ( .IN1(n825), .IN2(C1_DATA9_0), .IN3(n509), .OUT(n510) );
  NAND3X1 U913 ( .IN1(n515), .IN2(n514), .IN3(n513), .OUT(n516) );
  AOI21 U914 ( .IN1(n835), .IN2(C1_DATA9_0), .IN3(n516), .OUT(n525) );
  INVX4 U915 ( .IN(n619), .OUT(n842) );
  AOI22 U916 ( .IN1(n916), .IN2(Datain1[7]), .IN3(Datain2[7]), .IN4(n957), 
        .OUT(n522) );
  AOI21 U917 ( .IN1(N360), .IN2(n842), .IN3(n523), .OUT(n524) );
  OAI21 U918 ( .IN1(n653), .IN2(n525), .IN3(n524), .OUT(n547) );
  OAI21 U919 ( .IN1(n179), .IN2(n180), .IN3(n526), .OUT(n527) );
  AOI22 U920 ( .IN1(n988), .IN2(n530), .IN3(n987), .IN4(n529), .OUT(n531) );
  INVX4 U921 ( .IN(Multi_ack), .OUT(n1015) );
  OAI21 U922 ( .IN1(n752), .IN2(n921), .IN3(n844), .OUT(n544) );
  NAND3X1 U923 ( .IN1(n536), .IN2(n705), .IN3(n676), .OUT(n537) );
  NAND3X1 U924 ( .IN1(n538), .IN2(n700), .IN3(n681), .OUT(n539) );
  INVX4 U925 ( .IN(n569), .OUT(n781) );
  MUX2X1 U926 ( .IN1(n816), .IN2(n781), .S(C1_DATA9_0), .OUT(n546) );
  NOR2X1 U927 ( .IN1(n547), .IN2(n546), .OUT(n553) );
  NAND3X1 U928 ( .IN1(n845), .IN2(n850), .IN3(n841), .OUT(n552) );
  AOI21 U929 ( .IN1(n781), .IN2(DP_OP_345_166_2358_n31), .IN3(n816), .OUT(n635) );
  AOI22 U930 ( .IN1(n832), .IN2(C1_DATA2_1), .IN3(n831), .IN4(C1_DATA2_1), 
        .OUT(n562) );
  AOI22 U931 ( .IN1(n834), .IN2(n404), .IN3(n404), .IN4(n833), .OUT(n559) );
  AOI22 U932 ( .IN1(n820), .IN2(C1_DATA1_1), .IN3(C1_DATA2_1), .IN4(n822), 
        .OUT(n556) );
  AOI22 U933 ( .IN1(n821), .IN2(C1_DATA5_1), .IN3(n817), .IN4(n404), .OUT(n554) );
  NAND3X1 U934 ( .IN1(n556), .IN2(n555), .IN3(n554), .OUT(n557) );
  AOI21 U935 ( .IN1(n825), .IN2(C1_DATA11_1), .IN3(n557), .OUT(n558) );
  NAND3X1 U936 ( .IN1(n563), .IN2(n562), .IN3(n561), .OUT(n564) );
  AOI21 U937 ( .IN1(n835), .IN2(C1_DATA13_1), .IN3(n564), .OUT(n566) );
  OAI21 U938 ( .IN1(n653), .IN2(n566), .IN3(n565), .OUT(n567) );
  NOR2X1 U939 ( .IN1(n567), .IN2(n654), .OUT(n568) );
  OAI21 U940 ( .IN1(n635), .IN2(n190), .IN3(n568), .OUT(n692) );
  AOI22 U941 ( .IN1(n916), .IN2(Datain1[12]), .IN3(Datain2[12]), .IN4(n957), 
        .OUT(n582) );
  NOR2X1 U942 ( .IN1(n782), .IN2(n569), .OUT(n584) );
  NAND3X1 U943 ( .IN1(n599), .IN2(DP_OP_349_170_2358_n56), .IN3(n584), .OUT(
        n581) );
  AOI22 U944 ( .IN1(n820), .IN2(C1_DATA1_5), .IN3(C1_DATA5_5), .IN4(n821), 
        .OUT(n570) );
  AOI21 U945 ( .IN1(n825), .IN2(C1_DATA11_5), .IN3(n571), .OUT(n573) );
  AOI22 U946 ( .IN1(n827), .IN2(C1_DATA7_5), .IN3(n826), .IN4(C1_DATA9_5), 
        .OUT(n572) );
  NAND3X1 U947 ( .IN1(n574), .IN2(n573), .IN3(n572), .OUT(n579) );
  AOI22 U948 ( .IN1(n832), .IN2(C1_DATA6_5), .IN3(n831), .IN4(C1_DATA10_5), 
        .OUT(n577) );
  NAND3X1 U949 ( .IN1(n577), .IN2(n576), .IN3(n575), .OUT(n578) );
  INVX4 U950 ( .IN(n653), .OUT(n951) );
  OAI21 U951 ( .IN1(n579), .IN2(n578), .IN3(n951), .OUT(n580) );
  NAND3X1 U952 ( .IN1(n582), .IN2(n581), .IN3(n580), .OUT(n583) );
  AOI21 U953 ( .IN1(n842), .IN2(N365), .IN3(n583), .OUT(n586) );
  NAND3X1 U954 ( .IN1(n586), .IN2(n585), .IN3(n785), .OUT(n696) );
  AOI22 U955 ( .IN1(n834), .IN2(C1_DATA12_4), .IN3(C1_DATA8_4), .IN4(n833), 
        .OUT(n588) );
  AOI22 U956 ( .IN1(n832), .IN2(C1_DATA6_4), .IN3(n831), .IN4(C1_DATA10_4), 
        .OUT(n587) );
  AOI21 U957 ( .IN1(n835), .IN2(C1_DATA13_4), .IN3(n589), .OUT(n596) );
  AOI22 U958 ( .IN1(n822), .IN2(C1_DATA2_4), .IN3(C1_DATA4_4), .IN4(n817), 
        .OUT(n592) );
  AOI22 U959 ( .IN1(n827), .IN2(C1_DATA7_4), .IN3(n826), .IN4(C1_DATA9_4), 
        .OUT(n590) );
  NAND3X1 U960 ( .IN1(n592), .IN2(n591), .IN3(n590), .OUT(n593) );
  NOR2X1 U961 ( .IN1(n594), .IN2(n593), .OUT(n595) );
  AOI21 U962 ( .IN1(n596), .IN2(n595), .IN3(n653), .OUT(n597) );
  NOR2X1 U963 ( .IN1(n598), .IN2(n597), .OUT(n602) );
  AOI21 U964 ( .IN1(n781), .IN2(n649), .IN3(n816), .OUT(n657) );
  MUX2X1 U965 ( .IN1(n600), .IN2(n657), .S(DP_OP_349_170_2358_n56), .OUT(n601)
         );
  NAND3X1 U966 ( .IN1(n602), .IN2(n601), .IN3(n785), .OUT(n695) );
  AOI22 U967 ( .IN1(n916), .IN2(Datain1[14]), .IN3(n957), .IN4(Datain2[14]), 
        .OUT(n618) );
  OAI21 U968 ( .IN1(n184), .IN2(n603), .IN3(n178), .OUT(n604) );
  NAND3X1 U969 ( .IN1(n605), .IN2(n604), .IN3(n781), .OUT(n617) );
  AOI22 U970 ( .IN1(n818), .IN2(C1_DATA3_7), .IN3(C1_DATA4_7), .IN4(n817), 
        .OUT(n606) );
  AOI21 U971 ( .IN1(n821), .IN2(C1_DATA5_7), .IN3(n607), .OUT(n611) );
  AOI21 U972 ( .IN1(n825), .IN2(C1_DATA11_7), .IN3(n608), .OUT(n610) );
  AOI22 U973 ( .IN1(n827), .IN2(C1_DATA7_7), .IN3(n826), .IN4(C1_DATA9_7), 
        .OUT(n609) );
  NAND3X1 U974 ( .IN1(n611), .IN2(n610), .IN3(n609), .OUT(n616) );
  AOI22 U975 ( .IN1(n832), .IN2(C1_DATA6_7), .IN3(n831), .IN4(C1_DATA10_7), 
        .OUT(n614) );
  AOI22 U976 ( .IN1(n834), .IN2(C1_DATA12_7), .IN3(C1_DATA8_7), .IN4(n833), 
        .OUT(n613) );
  NAND3X1 U977 ( .IN1(n614), .IN2(n613), .IN3(n612), .OUT(n615) );
  AOI22 U978 ( .IN1(n827), .IN2(C1_DATA7_2), .IN3(n826), .IN4(C1_DATA9_2), 
        .OUT(n629) );
  AOI22 U979 ( .IN1(n832), .IN2(C1_DATA6_2), .IN3(n831), .IN4(C1_DATA10_2), 
        .OUT(n628) );
  AOI22 U980 ( .IN1(n834), .IN2(n166), .IN3(n394), .IN4(n833), .OUT(n625) );
  AOI22 U981 ( .IN1(n820), .IN2(C1_DATA1_2), .IN3(C1_DATA2_2), .IN4(n822), 
        .OUT(n622) );
  AOI22 U982 ( .IN1(n821), .IN2(C1_DATA5_2), .IN3(n817), .IN4(n166), .OUT(n620) );
  NAND3X1 U983 ( .IN1(n622), .IN2(n621), .IN3(n620), .OUT(n623) );
  AOI21 U984 ( .IN1(n825), .IN2(C1_DATA11_2), .IN3(n623), .OUT(n624) );
  NAND3X1 U985 ( .IN1(n629), .IN2(n628), .IN3(n627), .OUT(n630) );
  AOI21 U986 ( .IN1(n835), .IN2(C1_DATA13_2), .IN3(n630), .OUT(n631) );
  NOR2X1 U987 ( .IN1(n653), .IN2(n631), .OUT(n632) );
  NOR2X1 U988 ( .IN1(n633), .IN2(n632), .OUT(n637) );
  MUX2X1 U989 ( .IN1(n635), .IN2(n634), .S(n406), .OUT(n636) );
  NAND3X1 U990 ( .IN1(n637), .IN2(n636), .IN3(n785), .OUT(n693) );
  AOI22 U991 ( .IN1(n827), .IN2(C1_DATA7_3), .IN3(n826), .IN4(C1_DATA9_3), 
        .OUT(n647) );
  AOI22 U992 ( .IN1(n834), .IN2(C1_DATA12_3), .IN3(n165), .IN4(n833), .OUT(
        n643) );
  AOI22 U993 ( .IN1(n820), .IN2(C1_DATA1_3), .IN3(C1_DATA2_3), .IN4(n822), 
        .OUT(n640) );
  AOI22 U994 ( .IN1(n821), .IN2(C1_DATA5_3), .IN3(n817), .IN4(C1_DATA4_3), 
        .OUT(n638) );
  NAND3X1 U995 ( .IN1(n640), .IN2(n639), .IN3(n638), .OUT(n641) );
  AOI21 U996 ( .IN1(n825), .IN2(C1_DATA11_3), .IN3(n641), .OUT(n642) );
  NAND3X1 U997 ( .IN1(n647), .IN2(n646), .IN3(n645), .OUT(n648) );
  AOI21 U998 ( .IN1(n835), .IN2(C1_DATA13_3), .IN3(n648), .OUT(n652) );
  OAI21 U999 ( .IN1(n653), .IN2(n652), .IN3(n651), .OUT(n655) );
  NOR2X1 U1000 ( .IN1(n655), .IN2(n654), .OUT(n656) );
  OAI21 U1001 ( .IN1(n657), .IN2(n407), .IN3(n656), .OUT(n694) );
  NAND3X1 U1002 ( .IN1(n658), .IN2(n728), .IN3(n711), .OUT(n671) );
  NOR2X1 U1003 ( .IN1(n672), .IN2(n671), .OUT(n673) );
  NOR2X1 U1004 ( .IN1(n678), .IN2(n677), .OUT(n680) );
  OAI21 U1005 ( .IN1(n701), .IN2(n700), .IN3(n681), .OUT(n703) );
  NOR2X1 U1006 ( .IN1(n703), .IN2(n702), .OUT(n704) );
  OAI21 U1007 ( .IN1(n706), .IN2(n705), .IN3(n704), .OUT(n707) );
  NAND3X1 U1008 ( .IN1(n714), .IN2(n713), .IN3(n712), .OUT(n715) );
  NOR2X1 U1009 ( .IN1(n716), .IN2(n715), .OUT(n717) );
  NAND3X1 U1010 ( .IN1(n720), .IN2(n718), .IN3(n719), .OUT(n727) );
  AOI21 U1011 ( .IN1(n396), .IN2(n723), .IN3(n722), .OUT(n726) );
  NOR2X1 U1012 ( .IN1(n930), .IN2(n861), .OUT(n730) );
  NOR2X1 U1013 ( .IN1(n734), .IN2(n869), .OUT(n739) );
  AOI22 U1014 ( .IN1(n403), .IN2(n848), .IN3(Multi_dataout[6]), .IN4(n894), 
        .OUT(n736) );
  AOI21 U1015 ( .IN1(n913), .IN2(n946), .IN3(n737), .OUT(n742) );
  AOI21 U1016 ( .IN1(n738), .IN2(n1014), .IN3(RSTn_BAR), .OUT(n749) );
  INVX4 U1017 ( .IN(n911), .OUT(n945) );
  AOI22 U1018 ( .IN1(G_reg), .IN2(n749), .IN3(n171), .IN4(n912), .OUT(n741) );
  OAI21 U1019 ( .IN1(RSTn_BAR), .IN2(n742), .IN3(n741), .OUT(n97) );
  AOI22 U1020 ( .IN1(Multi_dataout[6]), .IN2(n848), .IN3(n391), .IN4(n894), 
        .OUT(n745) );
  OAI21 U1021 ( .IN1(n746), .IN2(n948), .IN3(n745), .OUT(n747) );
  NAND3X1 U1022 ( .IN1(n801), .IN2(n200), .IN3(n788), .OUT(n764) );
  NAND3X1 U1023 ( .IN1(Multi_ack), .IN2(Multi_dataout[15]), .IN3(n751), .OUT(
        n750) );
  NAND3X1 U1024 ( .IN1(n754), .IN2(n753), .IN3(n759), .OUT(n795) );
  AOI21 U1025 ( .IN1(n791), .IN2(Exc_value[0]), .IN3(n756), .OUT(n761) );
  NAND3X1 U1026 ( .IN1(n761), .IN2(n799), .IN3(n792), .OUT(n762) );
  AOI21 U1027 ( .IN1(n200), .IN2(n795), .IN3(n762), .OUT(n763) );
  AOI21 U1028 ( .IN1(n764), .IN2(n763), .IN3(RSTn_BAR), .OUT(n765) );
  AOI22 U1029 ( .IN1(n916), .IN2(Datain1[13]), .IN3(n957), .IN4(Datain2[13]), 
        .OUT(n779) );
  AOI22 U1030 ( .IN1(n818), .IN2(C1_DATA3_6), .IN3(C1_DATA4_6), .IN4(n817), 
        .OUT(n766) );
  AOI21 U1031 ( .IN1(n821), .IN2(C1_DATA5_6), .IN3(n767), .OUT(n772) );
  AOI21 U1032 ( .IN1(n825), .IN2(C1_DATA11_6), .IN3(n769), .OUT(n771) );
  AOI22 U1033 ( .IN1(n827), .IN2(C1_DATA7_6), .IN3(n826), .IN4(C1_DATA9_6), 
        .OUT(n770) );
  NAND3X1 U1034 ( .IN1(n772), .IN2(n771), .IN3(n770), .OUT(n777) );
  AOI22 U1035 ( .IN1(n832), .IN2(C1_DATA6_6), .IN3(n831), .IN4(C1_DATA10_6), 
        .OUT(n775) );
  AOI22 U1036 ( .IN1(n834), .IN2(C1_DATA12_6), .IN3(C1_DATA8_6), .IN4(n833), 
        .OUT(n774) );
  NAND3X1 U1037 ( .IN1(n775), .IN2(n774), .IN3(n773), .OUT(n776) );
  OAI21 U1038 ( .IN1(n776), .IN2(n777), .IN3(n951), .OUT(n778) );
  AOI21 U1039 ( .IN1(n842), .IN2(N366), .IN3(n780), .OUT(n787) );
  MUX2X1 U1040 ( .IN1(n784), .IN2(n783), .S(DP_OP_349_170_2358_n58), .OUT(n786) );
  NAND3X1 U1041 ( .IN1(n787), .IN2(n786), .IN3(n785), .OUT(n697) );
  NAND3X1 U1042 ( .IN1(n789), .IN2(n193), .IN3(n788), .OUT(n797) );
  AOI21 U1043 ( .IN1(n791), .IN2(Exc_value[2]), .IN3(n790), .OUT(n793) );
  AOI21 U1044 ( .IN1(n795), .IN2(n193), .IN3(n794), .OUT(n796) );
  AOI21 U1045 ( .IN1(n797), .IN2(n796), .IN3(RSTn_BAR), .OUT(n798) );
  NAND3X1 U1046 ( .IN1(n921), .IN2(n990), .IN3(n799), .OUT(n800) );
  AOI21 U1047 ( .IN1(N368), .IN2(n801), .IN3(n800), .OUT(n815) );
  NAND3X1 U1048 ( .IN1(n206), .IN2(n205), .IN3(n203), .OUT(n802) );
  AOI21 U1049 ( .IN1(n803), .IN2(n802), .IN3(n1013), .OUT(n804) );
  OAI21 U1050 ( .IN1(n849), .IN2(n805), .IN3(n804), .OUT(n806) );
  NOR2X1 U1051 ( .IN1(n1030), .IN2(n806), .OUT(n807) );
  AOI21 U1052 ( .IN1(n815), .IN2(n807), .IN3(RSTn_BAR), .OUT(n808) );
  OAI21 U1053 ( .IN1(n809), .IN2(n1024), .IN3(n987), .OUT(n811) );
  NAND3X1 U1054 ( .IN1(n812), .IN2(n811), .IN3(n810), .OUT(n813) );
  AOI21 U1055 ( .IN1(n815), .IN2(n814), .IN3(RSTn_BAR), .OUT(N72) );
  AOI21 U1056 ( .IN1(n820), .IN2(C1_DATA1_8), .IN3(n819), .OUT(n830) );
  AOI22 U1057 ( .IN1(n822), .IN2(C1_DATA2_8), .IN3(C1_DATA5_8), .IN4(n821), 
        .OUT(n823) );
  AOI21 U1058 ( .IN1(n825), .IN2(C1_DATA11_8), .IN3(n824), .OUT(n829) );
  AOI22 U1059 ( .IN1(n827), .IN2(C1_DATA7_8), .IN3(n826), .IN4(C1_DATA9_8), 
        .OUT(n828) );
  NAND3X1 U1060 ( .IN1(n830), .IN2(n829), .IN3(n828), .OUT(n840) );
  AOI22 U1061 ( .IN1(n832), .IN2(C1_DATA6_8), .IN3(n831), .IN4(C1_DATA10_8), 
        .OUT(n838) );
  AOI22 U1062 ( .IN1(n834), .IN2(C1_DATA12_8), .IN3(C1_DATA8_8), .IN4(n833), 
        .OUT(n837) );
  NAND3X1 U1063 ( .IN1(n838), .IN2(n837), .IN3(n836), .OUT(n839) );
  NAND3X1 U1064 ( .IN1(G_reg), .IN2(T_reg), .IN3(n401), .OUT(n847) );
  AOI21 U1065 ( .IN1(n401), .IN2(n188), .IN3(n878), .OUT(n846) );
  MUX2X1 U1066 ( .IN1(n847), .IN2(n846), .S(Final_Mantissa_reg[0]), .OUT(n857)
         );
  OAI21 U1067 ( .IN1(n851), .IN2(n936), .IN3(n850), .OUT(n852) );
  AOI21 U1068 ( .IN1(Datain2[0]), .IN2(n938), .IN3(n852), .OUT(n853) );
  OAI21 U1069 ( .IN1(n854), .IN2(n910), .IN3(n853), .OUT(n855) );
  AOI21 U1070 ( .IN1(n922), .IN2(Multi_dataout[8]), .IN3(n855), .OUT(n856) );
  AOI21 U1071 ( .IN1(G_reg), .IN2(Final_Mantissa_reg[0]), .IN3(
        Final_Mantissa_reg[1]), .OUT(n859) );
  NOR2X1 U1072 ( .IN1(n859), .IN2(n890), .OUT(n860) );
  AOI22 U1073 ( .IN1(n401), .IN2(n860), .IN3(Multi_dataout[8]), .IN4(n894), 
        .OUT(n876) );
  NOR2X1 U1074 ( .IN1(n862), .IN2(n861), .OUT(n867) );
  OAI21 U1075 ( .IN1(n865), .IN2(n864), .IN3(DP_OP_349_170_2358_n55), .OUT(
        n866) );
  AOI21 U1076 ( .IN1(n941), .IN2(n946), .IN3(n877), .OUT(n885) );
  AOI22 U1077 ( .IN1(n916), .IN2(Datain1[1]), .IN3(n957), .IN4(Datain2[1]), 
        .OUT(n881) );
  OAI21 U1078 ( .IN1(n199), .IN2(n882), .IN3(n881), .OUT(n883) );
  AOI21 U1079 ( .IN1(n397), .IN2(n171), .IN3(n883), .OUT(n884) );
  OAI21 U1080 ( .IN1(RSTn_BAR), .IN2(n885), .IN3(n884), .OUT(n686) );
  OAI21 U1081 ( .IN1(n890), .IN2(Final_Mantissa_reg[2]), .IN3(n907), .OUT(n892) );
  OAI21 U1082 ( .IN1(n892), .IN2(n952), .IN3(n891), .OUT(n893) );
  AOI21 U1083 ( .IN1(n957), .IN2(Datain2[2]), .IN3(n893), .OUT(n897) );
  NAND3X1 U1084 ( .IN1(n395), .IN2(n409), .IN3(n894), .OUT(n896) );
  NAND3X1 U1085 ( .IN1(Multi_dataout[10]), .IN2(n409), .IN3(n922), .OUT(n895)
         );
  NAND3X1 U1086 ( .IN1(n897), .IN2(n896), .IN3(n895), .OUT(n898) );
  AOI21 U1087 ( .IN1(Final_Mantissa_reg[2]), .IN2(n959), .IN3(n898), .OUT(n899) );
  AOI21 U1088 ( .IN1(n963), .IN2(n171), .IN3(n901), .OUT(n902) );
  OAI21 U1089 ( .IN1(n301), .IN2(n949), .IN3(n902), .OUT(n687) );
  AOI21 U1090 ( .IN1(n904), .IN2(n933), .IN3(n959), .OUT(n918) );
  AOI22 U1091 ( .IN1(n916), .IN2(Datain1[3]), .IN3(n957), .IN4(Datain2[3]), 
        .OUT(n905) );
  OAI21 U1092 ( .IN1(n195), .IN2(n918), .IN3(n905), .OUT(n906) );
  NOR2X1 U1093 ( .IN1(n924), .IN2(n921), .OUT(n908) );
  AOI22 U1094 ( .IN1(n909), .IN2(n908), .IN3(Multi_dataout[11]), .IN4(n922), 
        .OUT(n914) );
  AOI22 U1095 ( .IN1(n916), .IN2(Datain1[4]), .IN3(n957), .IN4(Datain2[4]), 
        .OUT(n917) );
  OAI21 U1096 ( .IN1(n187), .IN2(n918), .IN3(n917), .OUT(n919) );
  AOI21 U1097 ( .IN1(n171), .IN2(n920), .IN3(n919), .OUT(n929) );
  NOR2X1 U1098 ( .IN1(Final_Mantissa_reg[4]), .IN2(n921), .OUT(n923) );
  AOI22 U1099 ( .IN1(n924), .IN2(n923), .IN3(n159), .IN4(n922), .OUT(n927) );
  NOR2X1 U1100 ( .IN1(n931), .IN2(n930), .OUT(n932) );
  OAI21 U1101 ( .IN1(n187), .IN2(n933), .IN3(n197), .OUT(n934) );
  NAND3X1 U1102 ( .IN1(n401), .IN2(n934), .IN3(n953), .OUT(n935) );
  AOI21 U1103 ( .IN1(n198), .IN2(n953), .IN3(n952), .OUT(n955) );
  OAI21 U1104 ( .IN1(n968), .IN2(n967), .IN3(n402), .OUT(n969) );
  OAI21 U1105 ( .IN1(n204), .IN2(n970), .IN3(n969), .OUT(n685) );
  AOI22 U1106 ( .IN1(n402), .IN2(n971), .IN3(Op1_Mantissa_reg[7]), .IN4(n1009), 
        .OUT(n972) );
  AOI22 U1107 ( .IN1(n988), .IN2(Datain1[0]), .IN3(n987), .IN4(Datain2[0]), 
        .OUT(n973) );
  OAI21 U1108 ( .IN1(n196), .IN2(n990), .IN3(n973), .OUT(ExcCheck_Datain[0])
         );
  AOI22 U1109 ( .IN1(n988), .IN2(Datain1[1]), .IN3(n987), .IN4(Datain2[1]), 
        .OUT(n974) );
  OAI21 U1110 ( .IN1(n199), .IN2(n990), .IN3(n974), .OUT(ExcCheck_Datain[1])
         );
  AOI22 U1111 ( .IN1(n988), .IN2(Datain1[2]), .IN3(n987), .IN4(Datain2[2]), 
        .OUT(n975) );
  OAI21 U1112 ( .IN1(n194), .IN2(n990), .IN3(n975), .OUT(ExcCheck_Datain[2])
         );
  AOI22 U1113 ( .IN1(n988), .IN2(Datain1[3]), .IN3(n987), .IN4(Datain2[3]), 
        .OUT(n976) );
  OAI21 U1114 ( .IN1(n195), .IN2(n990), .IN3(n976), .OUT(ExcCheck_Datain[3])
         );
  AOI22 U1115 ( .IN1(n988), .IN2(Datain1[4]), .IN3(n987), .IN4(Datain2[4]), 
        .OUT(n977) );
  OAI21 U1116 ( .IN1(n187), .IN2(n990), .IN3(n977), .OUT(ExcCheck_Datain[4])
         );
  AOI22 U1117 ( .IN1(n988), .IN2(Datain1[5]), .IN3(n987), .IN4(Datain2[5]), 
        .OUT(n978) );
  OAI21 U1118 ( .IN1(n197), .IN2(n990), .IN3(n978), .OUT(ExcCheck_Datain[5])
         );
  AOI22 U1119 ( .IN1(n988), .IN2(Datain1[6]), .IN3(n987), .IN4(Datain2[6]), 
        .OUT(n979) );
  OAI21 U1120 ( .IN1(n198), .IN2(n990), .IN3(n979), .OUT(ExcCheck_Datain[6])
         );
  AOI22 U1121 ( .IN1(n988), .IN2(Datain1[7]), .IN3(Datain2[7]), .IN4(n987), 
        .OUT(n980) );
  OAI21 U1122 ( .IN1(C1_DATA9_0), .IN2(n990), .IN3(n980), .OUT(
        ExcCheck_Datain[7]) );
  AOI22 U1123 ( .IN1(n987), .IN2(Datain2[8]), .IN3(Datain1[8]), .IN4(n988), 
        .OUT(n981) );
  OAI21 U1124 ( .IN1(C1_DATA2_1), .IN2(n990), .IN3(n981), .OUT(
        ExcCheck_Datain[8]) );
  AOI22 U1125 ( .IN1(n987), .IN2(Datain2[9]), .IN3(Datain1[9]), .IN4(n988), 
        .OUT(n982) );
  OAI21 U1126 ( .IN1(n406), .IN2(n990), .IN3(n982), .OUT(ExcCheck_Datain[9])
         );
  AOI22 U1127 ( .IN1(n988), .IN2(Datain1[10]), .IN3(n987), .IN4(Datain2[10]), 
        .OUT(n983) );
  OAI21 U1128 ( .IN1(n407), .IN2(n990), .IN3(n983), .OUT(ExcCheck_Datain[10])
         );
  AOI22 U1129 ( .IN1(n988), .IN2(Datain1[11]), .IN3(n987), .IN4(Datain2[11]), 
        .OUT(n984) );
  OAI21 U1130 ( .IN1(n183), .IN2(n990), .IN3(n984), .OUT(ExcCheck_Datain[11])
         );
  AOI22 U1131 ( .IN1(n988), .IN2(Datain1[12]), .IN3(Datain2[12]), .IN4(n987), 
        .OUT(n985) );
  OAI21 U1132 ( .IN1(n185), .IN2(n990), .IN3(n985), .OUT(ExcCheck_Datain[12])
         );
  AOI22 U1133 ( .IN1(n988), .IN2(Datain1[13]), .IN3(n987), .IN4(Datain2[13]), 
        .OUT(n986) );
  OAI21 U1134 ( .IN1(n184), .IN2(n990), .IN3(n986), .OUT(ExcCheck_Datain[13])
         );
  AOI22 U1135 ( .IN1(n988), .IN2(Datain1[14]), .IN3(n987), .IN4(Datain2[14]), 
        .OUT(n989) );
  OAI21 U1136 ( .IN1(n178), .IN2(n990), .IN3(n989), .OUT(ExcCheck_Datain[14])
         );
  NOR2X1 U1137 ( .IN1(n1016), .IN2(Exc_value[1]), .OUT(n1017) );
  NAND2X1 U1138 ( .IN1(Datain1[10]), .IN2(Datain1[9]), .OUT(n1019) );
  NAND3X1 U1139 ( .IN1(Datain1[8]), .IN2(Datain1[13]), .IN3(Datain1[11]), 
        .OUT(n1018) );
  NOR2X1 U1140 ( .IN1(n1019), .IN2(n1018), .OUT(n1020) );
  NAND2X1 U1141 ( .IN1(Datain2[10]), .IN2(Datain2[11]), .OUT(n1022) );
  NAND3X1 U1142 ( .IN1(Datain2[13]), .IN2(Datain2[8]), .IN3(Datain2[9]), .OUT(
        n1021) );
  NOR2X1 U1143 ( .IN1(n1022), .IN2(n1021), .OUT(n1023) );
  AOI22 U1144 ( .IN1(n1025), .IN2(n401), .IN3(n1013), .IN4(n1024), .OUT(n1027)
         );
  AOI21 U1145 ( .IN1(Exc_Ack), .IN2(n1010), .IN3(n1012), .OUT(n1026) );
  NAND3X1 U1146 ( .IN1(n1027), .IN2(n1034), .IN3(n1026), .OUT(n1028) );
  NOR2X1 U1147 ( .IN1(n1028), .IN2(n1030), .OUT(n1029) );
  NOR2X1 U1148 ( .IN1(RSTn_BAR), .IN2(n1029), .OUT(N70) );
  NOR2X1 U1149 ( .IN1(n215), .IN2(n1031), .OUT(Dataout[15]) );
  AOI21 U1150 ( .IN1(n401), .IN2(n1032), .IN3(n1012), .OUT(n1033) );
  NOR2X1 U1151 ( .IN1(RSTn_BAR), .IN2(n1009), .OUT(n1059) );
  NOR2X1 U1152 ( .IN1(RSTn_BAR), .IN2(Exc_Ack), .OUT(n1039) );
  NAND3X1 U1153 ( .IN1(n1040), .IN2(n1036), .IN3(n1035), .OUT(n1037) );
  MUX2X1 U1154 ( .IN1(ExcCheck_valid), .IN2(n1039), .S(n1038), .OUT(n684) );
  OAI21 U1155 ( .IN1(Datain1[15]), .IN2(Datain2[15]), .IN3(n1040), .OUT(n1041)
         );
  AOI21 U1156 ( .IN1(Datain1[15]), .IN2(Datain2[15]), .IN3(n1041), .OUT(n1042)
         );
  NAND3X1 U1157 ( .IN1(n1014), .IN2(Data_valid), .IN3(n1042), .OUT(n1045) );
  AOI21 U1158 ( .IN1(n1045), .IN2(n1044), .IN3(RSTn_BAR), .OUT(n683) );
  NAND3X1 U1159 ( .IN1(n1062), .IN2(n409), .IN3(n1015), .OUT(n1061) );
  OAI21 U1160 ( .IN1(n1062), .IN2(n216), .IN3(n1061), .OUT(n682) );
  AOI22 U1161 ( .IN1(Datain2[6]), .IN2(n402), .IN3(Op2_Mantissa_reg[6]), .IN4(
        n1009), .OUT(n1046) );
  AOI22 U1162 ( .IN1(Datain2[5]), .IN2(n402), .IN3(Op2_Mantissa_reg[5]), .IN4(
        n1009), .OUT(n1047) );
  AOI22 U1163 ( .IN1(Datain2[4]), .IN2(n402), .IN3(Op2_Mantissa_reg[4]), .IN4(
        n1009), .OUT(n1048) );
  AOI22 U1164 ( .IN1(Datain2[3]), .IN2(n402), .IN3(Op2_Mantissa_reg[3]), .IN4(
        n1009), .OUT(n1049) );
  AOI22 U1165 ( .IN1(Datain2[2]), .IN2(n402), .IN3(Op2_Mantissa_reg[2]), .IN4(
        n1009), .OUT(n1050) );
  AOI22 U1166 ( .IN1(Datain2[1]), .IN2(n402), .IN3(Op2_Mantissa_reg[1]), .IN4(
        n1009), .OUT(n1051) );
  AOI22 U1167 ( .IN1(Datain2[0]), .IN2(n402), .IN3(Op2_Mantissa_reg[0]), .IN4(
        n1009), .OUT(n1052) );
  AOI22 U1168 ( .IN1(Datain1[6]), .IN2(n402), .IN3(Op1_Mantissa_reg[6]), .IN4(
        n1009), .OUT(n1053) );
  AOI22 U1169 ( .IN1(Datain1[5]), .IN2(n402), .IN3(Op1_Mantissa_reg[5]), .IN4(
        n1009), .OUT(n1054) );
  AOI22 U1170 ( .IN1(Datain1[4]), .IN2(n402), .IN3(Op1_Mantissa_reg[4]), .IN4(
        n1009), .OUT(n1055) );
  AOI22 U1171 ( .IN1(Datain1[3]), .IN2(n402), .IN3(Op1_Mantissa_reg[3]), .IN4(
        n1009), .OUT(n1056) );
  AOI22 U1172 ( .IN1(Datain1[2]), .IN2(n402), .IN3(Op1_Mantissa_reg[2]), .IN4(
        n1009), .OUT(n1057) );
  AOI22 U1173 ( .IN1(Datain1[1]), .IN2(n402), .IN3(Op1_Mantissa_reg[1]), .IN4(
        n1009), .OUT(n1058) );
  AOI22 U1174 ( .IN1(Datain1[0]), .IN2(n402), .IN3(Op1_Mantissa_reg[0]), .IN4(
        n1009), .OUT(n1060) );
  OAI21 U1175 ( .IN1(RSTn_BAR), .IN2(n1015), .IN3(n1062), .OUT(n1078) );
  AOI22 U1176 ( .IN1(Op2_Mantissa_reg[7]), .IN2(n1079), .IN3(Multi_datain2[7]), 
        .IN4(n1078), .OUT(n1063) );
  AOI22 U1177 ( .IN1(Op2_Mantissa_reg[6]), .IN2(n1079), .IN3(Multi_datain2[6]), 
        .IN4(n1078), .OUT(n1064) );
  AOI22 U1178 ( .IN1(Op2_Mantissa_reg[5]), .IN2(n1079), .IN3(Multi_datain2[5]), 
        .IN4(n1078), .OUT(n1065) );
  AOI22 U1179 ( .IN1(Op2_Mantissa_reg[4]), .IN2(n1079), .IN3(Multi_datain2[4]), 
        .IN4(n1078), .OUT(n1066) );
  AOI22 U1180 ( .IN1(Op2_Mantissa_reg[3]), .IN2(n1079), .IN3(Multi_datain2[3]), 
        .IN4(n1078), .OUT(n1067) );
  AOI22 U1181 ( .IN1(Op2_Mantissa_reg[2]), .IN2(n1079), .IN3(Multi_datain2[2]), 
        .IN4(n1078), .OUT(n1068) );
  AOI22 U1182 ( .IN1(Op2_Mantissa_reg[1]), .IN2(n1079), .IN3(Multi_datain2[1]), 
        .IN4(n1078), .OUT(n1069) );
  AOI22 U1183 ( .IN1(Op2_Mantissa_reg[0]), .IN2(n1079), .IN3(Multi_datain2[0]), 
        .IN4(n1078), .OUT(n1070) );
  AOI22 U1184 ( .IN1(Op1_Mantissa_reg[7]), .IN2(n1079), .IN3(Multi_datain1[7]), 
        .IN4(n1078), .OUT(n1071) );
  AOI22 U1185 ( .IN1(Op1_Mantissa_reg[6]), .IN2(n1079), .IN3(Multi_datain1[6]), 
        .IN4(n1078), .OUT(n1072) );
  AOI22 U1186 ( .IN1(Op1_Mantissa_reg[5]), .IN2(n1079), .IN3(Multi_datain1[5]), 
        .IN4(n1078), .OUT(n1073) );
  AOI22 U1187 ( .IN1(Op1_Mantissa_reg[4]), .IN2(n1079), .IN3(Multi_datain1[4]), 
        .IN4(n1078), .OUT(n1074) );
  AOI22 U1188 ( .IN1(Op1_Mantissa_reg[3]), .IN2(n1079), .IN3(Multi_datain1[3]), 
        .IN4(n1078), .OUT(n1075) );
  AOI22 U1189 ( .IN1(Op1_Mantissa_reg[2]), .IN2(n1079), .IN3(Multi_datain1[2]), 
        .IN4(n1078), .OUT(n1076) );
  AOI22 U1190 ( .IN1(Op1_Mantissa_reg[1]), .IN2(n1079), .IN3(Multi_datain1[1]), 
        .IN4(n1078), .OUT(n1077) );
  AOI22 U1191 ( .IN1(Op1_Mantissa_reg[0]), .IN2(n1079), .IN3(Multi_datain1[0]), 
        .IN4(n1078), .OUT(n1080) );
endmodule


module FPU_Control ( CLK, RSTn, CS, DIN1, DIN2, DIV, DACK, DR, DOUT, DOV, DOA, 
        ABUSY, MBUSY, EXC, OPT, MODE, DEBUG );
  input [15:0] DIN1;
  input [15:0] DIN2;
  output [15:0] DOUT;
  output [2:0] EXC;
  input [2:0] MODE;
  output [4:0] DEBUG;
  input CLK, RSTn, CS, DIV, DOA, OPT;
  output DACK, DR, DOV, ABUSY, MBUSY;
  wire   Add_carryout, N147, N148, N149, N150, N189, N190, N191,
         MulCntrl_valid, AdderCntrl_valid, AdderCntrl_Dataout_valid,
         MulCntrl_Dataout_valid, Add_valid, Add_ack, AdderCntrl_ExcCheck_valid,
         AdderCntrl_Exc_Ack, Booth_valid, Booth_ack, MulCntrl_ExcCheck_valid,
         MulCntrl_Exc_Ack, ExcSelect, ExcCheck_valid, AddSelect,
         u_exc_check_N45, u_exc_check_StateMC_0_,
         u_ExcChecker_interconnect_N53, u_ExcChecker_interconnect_priority_reg,
         u_ExcChecker_interconnect_stateMC_0_,
         u_ExcChecker_interconnect_stateMC_1_, u_booth_N258, u_booth_N55,
         u_booth_N54, u_booth_N53, u_booth_N52, u_booth_N51, u_booth_N50,
         u_booth_N49, u_booth_BStateMC_1_, u_booth_count_reg_2_,
         u_booth_count_reg_3_, u_booth_Q1_reg, u_booth_M_reg_1_,
         u_booth_M_reg_2_, u_booth_M_reg_3_, u_booth_M_reg_4_,
         u_booth_M_reg_5_, u_booth_M_reg_6_, u_booth_M_reg_7_,
         u_booth_A_reg_7_, u_booth_A_reg_8_, u_adder_24b_N131,
         u_adder_24b_N129, u_adder_24b_N122, u_adder_24b_StateMC_1_,
         u_Adder_interconnect_N53, u_Adder_interconnect_priority_reg,
         u_Adder_interconnect_stateMC_1_, n408, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n462, n463, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n587, n588, n592, n594, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n609, n610, n611, n612, n613, n614, n615,
         n616, n622, n654, n692, n694, n695, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n709, n710, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n734, n768, n802, n806, n992, n1021, n1028, n1031, n1034, n1037,
         n1040, n1043, n1078, n1080, n1089, n1092, n1135, n1302, n1513, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1587, n1588, n1589, n1620, n1621, n1622, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1692, n1723,
         add_x_173_n71, add_x_173_n69, add_x_173_n65, add_x_173_n64,
         add_x_173_n63, add_x_173_n61, add_x_173_n60, add_x_173_n59,
         add_x_173_n58, add_x_173_n57, add_x_173_n56, add_x_173_n55,
         add_x_173_n52, add_x_173_n51, add_x_173_n49, add_x_173_n48,
         add_x_173_n44, add_x_173_n43, add_x_173_n42, add_x_173_n41,
         add_x_173_n40, add_x_173_n39, add_x_173_n37, add_x_173_n36,
         add_x_173_n35, add_x_173_n34, add_x_173_n33, add_x_173_n31,
         add_x_173_n30, add_x_173_n23, add_x_173_n1, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7;
  wire   [8:0] Add_dataout;
  wire   [4:0] AdderCntrl_Debug;
  wire   [1:0] multStateMC;
  wire   [15:0] AdderCntrl_Op1;
  wire   [15:0] AdderCntrl_Op2;
  wire   [15:0] MulCntrl_Op1;
  wire   [15:0] MulCntrl_Op2;
  wire   [1:0] getdataStat_reg;
  wire   [15:0] AdderResult_reg;
  wire   [15:0] MultResult_reg;
  wire   [2:0] AddExc_reg;
  wire   [2:0] MultExc_reg;
  wire   [15:0] AdderCntrl_Dataout;
  wire   [2:0] AdderCntrl_Exc;
  wire   [15:0] MulCntrl_Dataout;
  wire   [2:0] MulCntrl_Exc;
  wire   [7:0] Add_Op1;
  wire   [8:0] Add_Op2;
  wire   [14:0] AdderCntrl_ExcCheck_Datain;
  wire   [2:0] ExcCheck_value;
  wire   [7:0] Booth_datain1;
  wire   [7:0] Booth_datain2;
  wire   [15:0] Booth_dataout;
  wire   [14:0] MulCntrl_ExcCheck_Datain;
  wire   [8:0] Booth_Add_datain1;
  wire   [8:0] Booth_Add_datain2;
  wire   [8:0] Add_Op1_wire;
  wire   [8:0] Add_Op2_wire;

  Adder_cntrl u_adder_cntrl ( .CLK(CLK), .Datain1({AdderCntrl_Op1[15:10], 
        n1869, n1871, AdderCntrl_Op1[7:0]}), .Datain2({AdderCntrl_Op2[15:9], 
        n1870, AdderCntrl_Op2[7:0]}), .Data_valid(AdderCntrl_valid), .Dataout(
        AdderCntrl_Dataout), .Exc(AdderCntrl_Exc), .Mode(MODE), .Debug(
        AdderCntrl_Debug), .Adder_datain1({SYNOPSYS_UNCONNECTED_1, Add_Op1}), 
        .Adder_datain2(Add_Op2), .Adder_valid(Add_valid), .Adder_dataout(
        Add_dataout), .Adder_carryout(Add_carryout), .Adder_ack(Add_ack), 
        .ExcCheck_valid(AdderCntrl_ExcCheck_valid), .Exc_value(ExcCheck_value), 
        .Exc_Ack(AdderCntrl_Exc_Ack), .RSTn_BAR(n1877), .Dataout_valid_BAR(
        AdderCntrl_Dataout_valid), .ExcCheck_Datain_14_(
        AdderCntrl_ExcCheck_Datain[14]), .ExcCheck_Datain_13__BAR(
        AdderCntrl_ExcCheck_Datain[13]), .ExcCheck_Datain_12_(
        AdderCntrl_ExcCheck_Datain[12]), .ExcCheck_Datain_11_(
        AdderCntrl_ExcCheck_Datain[11]), .ExcCheck_Datain_9_(
        AdderCntrl_ExcCheck_Datain[9]), .ExcCheck_Datain_8_(
        AdderCntrl_ExcCheck_Datain[8]), .ExcCheck_Datain_6_(
        AdderCntrl_ExcCheck_Datain[6]), .ExcCheck_Datain_5_(
        AdderCntrl_ExcCheck_Datain[5]), .ExcCheck_Datain_4_(
        AdderCntrl_ExcCheck_Datain[4]), .ExcCheck_Datain_3_(
        AdderCntrl_ExcCheck_Datain[3]), .ExcCheck_Datain_2_(
        AdderCntrl_ExcCheck_Datain[2]), .ExcCheck_Datain_1_(
        AdderCntrl_ExcCheck_Datain[1]), .ExcCheck_Datain_0_(
        AdderCntrl_ExcCheck_Datain[0]), .ExcCheck_Datain_10__BAR(
        AdderCntrl_ExcCheck_Datain[10]), .ExcCheck_Datain_7__BAR(
        AdderCntrl_ExcCheck_Datain[7]) );
  Mul_cntrl u_mul_cntrl ( .CLK(CLK), .Datain1({MulCntrl_Op1[15:9], n1865, 
        MulCntrl_Op1[7:0]}), .Datain2({MulCntrl_Op2[15:14], n1863, 
        MulCntrl_Op2[12:9], n1862, MulCntrl_Op2[7:0]}), .Data_valid(
        MulCntrl_valid), .Dataout(MulCntrl_Dataout), .Dataout_valid(
        MulCntrl_Dataout_valid), .Exc(MulCntrl_Exc), .Mode({n2293, n2293, 
        n2293}), .Debug({SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6}), .Multi_datain1(Booth_datain1), .Multi_datain2(Booth_datain2), .Multi_valid(
        Booth_valid), .Multi_dataout({Booth_dataout[15:12], n1866, n1864, 
        Booth_dataout[9], n1867, Booth_dataout[7], n1868, Booth_dataout[5:0]}), 
        .Multi_ack(Booth_ack), .ExcCheck_valid(MulCntrl_ExcCheck_valid), 
        .ExcCheck_Datain({SYNOPSYS_UNCONNECTED_7, MulCntrl_ExcCheck_Datain}), 
        .Exc_value(ExcCheck_value), .Exc_Ack(MulCntrl_Exc_Ack), .RSTn_BAR(
        n1877) );
  DFFRX1 u_Adder_interconnect_M2_ack_reg ( .D(n1587), .CLK(CLK), .CLRB(n408), 
        .Q(n1846), .QB(n1808) );
  DFFRX1 u_booth_A_reg_reg_7_ ( .D(n1546), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_A_reg_7_), .QB(n1828) );
  DFFRX1 u_booth_A_reg_reg_6_ ( .D(n1547), .CLK(CLK), .CLRB(n408), .Q(n1851), 
        .QB(n729) );
  DFFRX1 u_booth_Q_reg_reg_7_ ( .D(n1021), .CLK(CLK), .CLRB(n408), .Q(n721), 
        .QB(n1830) );
  DFFRX1 u_booth_Q_reg_reg_6_ ( .D(n1028), .CLK(CLK), .CLRB(n408), .Q(n720), 
        .QB(n1831) );
  DFFRX1 u_booth_Q_reg_reg_5_ ( .D(n1031), .CLK(CLK), .CLRB(n408), .Q(n719), 
        .QB(n1832) );
  DFFRX1 u_booth_Q_reg_reg_4_ ( .D(n1034), .CLK(CLK), .CLRB(n408), .Q(n718), 
        .QB(n1833) );
  DFFRX1 u_booth_Q_reg_reg_3_ ( .D(n1037), .CLK(CLK), .CLRB(n408), .Q(n717), 
        .QB(n1834) );
  DFFRX1 u_booth_Q_reg_reg_2_ ( .D(n1040), .CLK(CLK), .CLRB(n408), .Q(n716), 
        .QB(n1835) );
  DFFRX1 u_booth_Q_reg_reg_1_ ( .D(n1043), .CLK(CLK), .CLRB(n408), .Q(n715), 
        .QB(n1836) );
  DFFRX1 u_booth_Q_reg_reg_0_ ( .D(n1135), .CLK(CLK), .CLRB(n408), .Q(n714), 
        .QB(n1806) );
  DFFRX1 u_booth_count_reg_reg_0_ ( .D(n1554), .CLK(CLK), .CLRB(n408), .QB(
        n694) );
  DFFRX1 u_booth_count_reg_reg_1_ ( .D(n1080), .CLK(CLK), .CLRB(n408), .Q(n695), .QB(n1790) );
  DFFRX1 u_booth_count_reg_reg_2_ ( .D(n1555), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_count_reg_2_) );
  DFFRX1 u_booth_count_reg_reg_3_ ( .D(n1092), .CLK(CLK), .CLRB(n408), .Q(
        n1840), .QB(u_booth_count_reg_3_) );
  DFFRX1 u_booth_BStateMC_reg_1_ ( .D(n1089), .CLK(CLK), .CLRB(n408), .Q(n1819), .QB(u_booth_BStateMC_1_) );
  DFFRX1 u_booth_BStateMC_reg_0_ ( .D(n1556), .CLK(CLK), .CLRB(n408), .Q(n1788), .QB(n734) );
  DFFRX1 u_booth_Q1_reg_reg ( .D(n1078), .CLK(CLK), .CLRB(n408), .Q(n1816), 
        .QB(u_booth_Q1_reg) );
  DFFRX1 u_booth_Adder_valid_reg ( .D(n1653), .CLK(CLK), .CLRB(n408), .Q(n1843), .QB(n692) );
  DFFRX1 u_Adder_interconnect_priority_reg_reg ( .D(n1620), .CLK(CLK), .CLRB(
        n408), .Q(u_Adder_interconnect_priority_reg), .QB(n1826) );
  DFFRX1 u_Adder_interconnect_stateMC_reg_0_ ( .D(n1621), .CLK(CLK), .CLRB(
        n408), .Q(n1809), .QB(n806) );
  DFFRX1 u_Adder_interconnect_M1_ack_reg ( .D(n594), .CLK(CLK), .CLRB(n408), 
        .Q(Add_ack) );
  DFFRX1 u_ExcChecker_interconnect_stateMC_reg_1_ ( .D(n1661), .CLK(CLK), 
        .CLRB(n408), .Q(u_ExcChecker_interconnect_stateMC_1_), .QB(n1827) );
  DFFRX1 u_ExcChecker_interconnect_priority_reg_reg ( .D(n1659), .CLK(CLK), 
        .CLRB(n408), .Q(u_ExcChecker_interconnect_priority_reg), .QB(n1825) );
  DFFRX1 u_ExcChecker_interconnect_stateMC_reg_0_ ( .D(n1660), .CLK(CLK), 
        .CLRB(n408), .Q(u_ExcChecker_interconnect_stateMC_0_), .QB(n1820) );
  DFFRX1 u_ExcChecker_interconnect_S_req_reg ( .D(
        u_ExcChecker_interconnect_N53), .CLK(CLK), .CLRB(n408), .Q(
        ExcCheck_valid) );
  DFFRX1 u_exc_check_ACK_reg ( .D(u_exc_check_N45), .CLK(CLK), .CLRB(n408), 
        .QB(n1823) );
  DFFRX1 u_ExcChecker_interconnect_M2_ack_reg ( .D(n1656), .CLK(CLK), .CLRB(
        n408), .Q(MulCntrl_Exc_Ack) );
  DFFRX1 u_exc_check_StateMC_reg_0_ ( .D(n622), .CLK(CLK), .CLRB(n408), .Q(
        u_exc_check_StateMC_0_), .QB(n1837) );
  DFFRX1 u_exc_check_StateMC_reg_1_ ( .D(n1657), .CLK(CLK), .CLRB(n408), .Q(
        n1850), .QB(n654) );
  DFFRX1 u_ExcChecker_interconnect_Select_reg ( .D(n1658), .CLK(CLK), .CLRB(
        n408), .Q(ExcSelect), .QB(n1821) );
  DFFRX1 u_exc_check_AEXC_reg_2_ ( .D(n588), .CLK(CLK), .CLRB(n408), .Q(
        ExcCheck_value[2]) );
  DFFRX1 u_exc_check_AEXC_reg_1_ ( .D(n1654), .CLK(CLK), .CLRB(n408), .Q(
        ExcCheck_value[1]), .QB(n1847) );
  DFFRX1 u_exc_check_AEXC_reg_0_ ( .D(n1655), .CLK(CLK), .CLRB(n408), .Q(
        ExcCheck_value[0]), .QB(n1824) );
  DFFRX1 u_ExcChecker_interconnect_M1_ack_reg ( .D(n592), .CLK(CLK), .CLRB(
        n408), .Q(AdderCntrl_Exc_Ack) );
  DFFRX1 u_Adder_interconnect_stateMC_reg_1_ ( .D(n1622), .CLK(CLK), .CLRB(
        n408), .Q(u_Adder_interconnect_stateMC_1_), .QB(n1822) );
  DFFRX1 u_Adder_interconnect_S_req_reg ( .D(u_Adder_interconnect_N53), .CLK(
        CLK), .CLRB(n408), .Q(n1813), .QB(n802) );
  DFFRX1 u_adder_24b_StateMC_reg_1_ ( .D(n1589), .CLK(CLK), .CLRB(n408), .Q(
        u_adder_24b_StateMC_1_) );
  DFFRX1 u_adder_24b_StateMC_reg_0_ ( .D(n1588), .CLK(CLK), .CLRB(n408), .Q(
        n1845), .QB(n768) );
  DFFRX1 u_adder_24b_ACK_reg ( .D(n2030), .CLK(CLK), .CLRB(n408), .QB(n1838)
         );
  DFFRX1 u_adder_24b_Z_reg_8_ ( .D(n598), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[8]) );
  DFFRX1 u_adder_24b_Z_reg_7_ ( .D(n599), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[7]) );
  DFFRX1 u_adder_24b_Z_reg_6_ ( .D(n600), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[6]) );
  DFFRX1 u_booth_A_reg_reg_5_ ( .D(n1548), .CLK(CLK), .CLRB(n408), .Q(n1810), 
        .QB(n728) );
  DFFRX1 u_booth_Adder_datain1_reg_5_ ( .D(u_booth_N54), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[5]) );
  DFFRX1 u_adder_24b_Z_reg_5_ ( .D(n601), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[5]) );
  DFFRX1 u_booth_A_reg_reg_4_ ( .D(n1549), .CLK(CLK), .CLRB(n408), .Q(n1842), 
        .QB(n727) );
  DFFRX1 u_booth_Adder_datain1_reg_4_ ( .D(u_booth_N53), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[4]) );
  DFFRX1 u_adder_24b_Z_reg_4_ ( .D(n602), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[4]) );
  DFFRX1 u_booth_A_reg_reg_3_ ( .D(n1550), .CLK(CLK), .CLRB(n408), .Q(n1811), 
        .QB(n726) );
  DFFRX1 u_booth_Adder_datain1_reg_3_ ( .D(u_booth_N52), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[3]) );
  DFFRX1 u_adder_24b_Z_reg_3_ ( .D(n603), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[3]) );
  DFFRX1 u_booth_A_reg_reg_2_ ( .D(n1551), .CLK(CLK), .CLRB(n408), .Q(n1839), 
        .QB(n725) );
  DFFRX1 u_booth_Adder_datain1_reg_2_ ( .D(u_booth_N51), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[2]) );
  DFFRX1 u_adder_24b_Z_reg_2_ ( .D(n604), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[2]) );
  DFFRX1 u_booth_A_reg_reg_1_ ( .D(n1552), .CLK(CLK), .CLRB(n408), .Q(n1812), 
        .QB(n724) );
  DFFRX1 u_booth_Adder_datain1_reg_1_ ( .D(u_booth_N50), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[1]) );
  DFFRX1 u_adder_24b_Z_reg_1_ ( .D(n605), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[1]) );
  DFFRX1 u_booth_A_reg_reg_0_ ( .D(n1553), .CLK(CLK), .CLRB(n408), .Q(n1841), 
        .QB(n723) );
  DFFRX1 u_booth_Adder_datain1_reg_0_ ( .D(u_booth_N49), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[0]) );
  DFFRX1 u_adder_24b_Z_reg_0_ ( .D(n596), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[0]) );
  DFFRX1 u_booth_Q_reg_reg_8_ ( .D(n1544), .CLK(CLK), .CLRB(n408), .Q(n1844), 
        .QB(n722) );
  DFFRX1 u_adder_24b_COUT_reg ( .D(n597), .CLK(CLK), .CLRB(n408), .Q(
        Add_carryout) );
  DFFRX1 outputRdy_reg_reg_0_ ( .D(N189), .CLK(CLK), .CLRB(n408), .QB(n587) );
  DFFRX1 getdataStat_reg_reg_0_ ( .D(N147), .CLK(CLK), .CLRB(n408), .Q(
        getdataStat_reg[0]) );
  DFFRX1 AdderCntrl_Op2_reg_0_ ( .D(n551), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[0]) );
  DFFRX1 AdderCntrl_Op2_reg_1_ ( .D(n550), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[1]) );
  DFFRX1 AdderCntrl_Op2_reg_2_ ( .D(n549), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[2]) );
  DFFRX1 AdderCntrl_Op2_reg_3_ ( .D(n548), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[3]) );
  DFFRX1 AdderCntrl_Op2_reg_4_ ( .D(n547), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[4]) );
  DFFRX1 AdderCntrl_Op2_reg_5_ ( .D(n546), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[5]) );
  DFFRX1 AdderCntrl_Op2_reg_6_ ( .D(n545), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[6]) );
  DFFRX1 AdderCntrl_Op2_reg_7_ ( .D(n544), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[7]) );
  DFFRX1 AdderCntrl_Op2_reg_8_ ( .D(n543), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[8]) );
  DFFRX1 AdderCntrl_Op2_reg_9_ ( .D(n542), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[9]) );
  DFFRX1 AdderCntrl_Op2_reg_10_ ( .D(n541), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[10]) );
  DFFRX1 AdderCntrl_Op2_reg_11_ ( .D(n540), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[11]) );
  DFFRX1 AdderCntrl_Op2_reg_12_ ( .D(n539), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[12]) );
  DFFRX1 AdderCntrl_Op2_reg_13_ ( .D(n538), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[13]) );
  DFFRX1 AdderCntrl_Op2_reg_14_ ( .D(n537), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[14]) );
  DFFRX1 AdderCntrl_Op2_reg_15_ ( .D(n536), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[15]) );
  DFFRX1 AdderCntrl_Op1_reg_0_ ( .D(n535), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[0]) );
  DFFRX1 AdderCntrl_Op1_reg_1_ ( .D(n534), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[1]) );
  DFFRX1 AdderCntrl_Op1_reg_2_ ( .D(n533), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[2]) );
  DFFRX1 AdderCntrl_Op1_reg_3_ ( .D(n532), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[3]) );
  DFFRX1 AdderCntrl_Op1_reg_4_ ( .D(n531), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[4]) );
  DFFRX1 AdderCntrl_Op1_reg_5_ ( .D(n530), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[5]) );
  DFFRX1 AdderCntrl_Op1_reg_6_ ( .D(n529), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[6]) );
  DFFRX1 AdderCntrl_Op1_reg_7_ ( .D(n528), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[7]) );
  DFFRX1 AdderCntrl_Op1_reg_8_ ( .D(n527), .CLK(CLK), .CLRB(n408), .QB(n1803)
         );
  DFFRX1 AdderCntrl_Op1_reg_9_ ( .D(n526), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[9]) );
  DFFRX1 AdderCntrl_Op1_reg_10_ ( .D(n525), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[10]) );
  DFFRX1 AdderCntrl_Op1_reg_11_ ( .D(n524), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[11]) );
  DFFRX1 AdderCntrl_Op1_reg_12_ ( .D(n523), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[12]) );
  DFFRX1 AdderCntrl_Op1_reg_13_ ( .D(n522), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[13]) );
  DFFRX1 AdderCntrl_Op1_reg_14_ ( .D(n521), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[14]) );
  DFFRX1 AdderCntrl_Op1_reg_15_ ( .D(n520), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[15]) );
  DFFRX1 ABUSY_reg ( .D(N149), .CLK(CLK), .CLRB(n408), .Q(ABUSY) );
  DFFRX1 adderStateMC_reg_0_ ( .D(n1302), .CLK(CLK), .CLRB(n408), .Q(n463) );
  DFFRX1 adderStateMC_reg_1_ ( .D(n1692), .CLK(CLK), .CLRB(n408), .Q(n1815), 
        .QB(n462) );
  DFFRX1 AddExc_reg_reg_2_ ( .D(n414), .CLK(CLK), .CLRB(n408), .Q(
        AddExc_reg[2]) );
  DFFRX1 AddExc_reg_reg_1_ ( .D(n413), .CLK(CLK), .CLRB(n408), .Q(
        AddExc_reg[1]) );
  DFFRX1 AddExc_reg_reg_0_ ( .D(n412), .CLK(CLK), .CLRB(n408), .Q(
        AddExc_reg[0]) );
  DFFRX1 AdderResult_reg_reg_0_ ( .D(n415), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[0]) );
  DFFRX1 AdderResult_reg_reg_1_ ( .D(n416), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[1]) );
  DFFRX1 AdderResult_reg_reg_2_ ( .D(n417), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[2]) );
  DFFRX1 AdderResult_reg_reg_3_ ( .D(n418), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[3]) );
  DFFRX1 AdderResult_reg_reg_4_ ( .D(n419), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[4]) );
  DFFRX1 AdderResult_reg_reg_5_ ( .D(n420), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[5]) );
  DFFRX1 AdderResult_reg_reg_6_ ( .D(n421), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[6]) );
  DFFRX1 AdderResult_reg_reg_7_ ( .D(n422), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[7]) );
  DFFRX1 AdderResult_reg_reg_8_ ( .D(n423), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[8]) );
  DFFRX1 AdderResult_reg_reg_9_ ( .D(n424), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[9]) );
  DFFRX1 AdderResult_reg_reg_10_ ( .D(n425), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[10]) );
  DFFRX1 AdderResult_reg_reg_11_ ( .D(n426), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[11]) );
  DFFRX1 AdderResult_reg_reg_12_ ( .D(n427), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[12]) );
  DFFRX1 AdderResult_reg_reg_13_ ( .D(n428), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[13]) );
  DFFRX1 AdderResult_reg_reg_14_ ( .D(n429), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[14]) );
  DFFRX1 AdderResult_reg_reg_15_ ( .D(n430), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[15]) );
  DFFRX1 u_booth_A_reg_reg_8_ ( .D(n1545), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_A_reg_8_), .QB(n1849) );
  DFFRX1 u_booth_Adder_datain2_reg_8_ ( .D(n705), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[8]) );
  DFFRX1 u_booth_M_reg_reg_0_ ( .D(n609), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_N258), .QB(n1814) );
  DFFRX1 u_booth_Adder_datain2_reg_0_ ( .D(n697), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[0]) );
  DFFRX1 u_booth_M_reg_reg_1_ ( .D(n610), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_1_), .QB(n1805) );
  DFFRX1 u_booth_Adder_datain2_reg_1_ ( .D(n698), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[1]) );
  DFFRX1 u_booth_M_reg_reg_2_ ( .D(n611), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_2_) );
  DFFRX1 u_booth_Adder_datain2_reg_2_ ( .D(n699), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[2]) );
  DFFRX1 u_booth_M_reg_reg_3_ ( .D(n612), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_3_) );
  DFFRX1 u_booth_Adder_datain2_reg_3_ ( .D(n700), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[3]) );
  DFFRX1 u_booth_M_reg_reg_4_ ( .D(n613), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_4_) );
  DFFRX1 u_booth_Adder_datain2_reg_4_ ( .D(n701), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[4]) );
  DFFRX1 u_booth_M_reg_reg_5_ ( .D(n614), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_5_) );
  DFFRX1 u_booth_Adder_datain2_reg_5_ ( .D(n702), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[5]) );
  DFFRX1 u_booth_M_reg_reg_6_ ( .D(n615), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_6_) );
  DFFRX1 u_booth_Adder_datain2_reg_6_ ( .D(n703), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[6]) );
  DFFRX1 u_booth_M_reg_reg_7_ ( .D(n616), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_7_), .QB(n1829) );
  DFFRX1 u_booth_Adder_datain2_reg_7_ ( .D(n704), .CLK(CLK), .CLRB(n408), .QB(
        n1818) );
  DFFRX1 multStateMC_reg_0_ ( .D(n992), .CLK(CLK), .CLRB(n408), .Q(n1817), 
        .QB(multStateMC[0]) );
  DFFRX1 outputRdy_reg_reg_1_ ( .D(N190), .CLK(CLK), .CLRB(n408), .Q(n1848), 
        .QB(n584) );
  DFFRX1 multStateMC_reg_1_ ( .D(n1513), .CLK(CLK), .CLRB(n408), .Q(
        multStateMC[1]), .QB(n1807) );
  DFFRX1 getdataStat_reg_reg_1_ ( .D(N148), .CLK(CLK), .CLRB(n408), .Q(
        getdataStat_reg[1]) );
  DFFRX1 MulCntrl_Op2_reg_0_ ( .D(n583), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[0]) );
  DFFRX1 MulCntrl_Op2_reg_1_ ( .D(n582), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[1]) );
  DFFRX1 MulCntrl_Op2_reg_2_ ( .D(n581), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[2]) );
  DFFRX1 MulCntrl_Op2_reg_3_ ( .D(n580), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[3]) );
  DFFRX1 MulCntrl_Op2_reg_4_ ( .D(n579), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[4]) );
  DFFRX1 MulCntrl_Op2_reg_5_ ( .D(n578), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[5]) );
  DFFRX1 MulCntrl_Op2_reg_6_ ( .D(n577), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[6]) );
  DFFRX1 MulCntrl_Op2_reg_7_ ( .D(n576), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[7]) );
  DFFRX1 MulCntrl_Op2_reg_8_ ( .D(n575), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[8]) );
  DFFRX1 MulCntrl_Op2_reg_9_ ( .D(n574), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[9]) );
  DFFRX1 MulCntrl_Op2_reg_10_ ( .D(n573), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[10]) );
  DFFRX1 MulCntrl_Op2_reg_11_ ( .D(n572), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[11]) );
  DFFRX1 MulCntrl_Op2_reg_12_ ( .D(n571), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[12]) );
  DFFRX1 MulCntrl_Op2_reg_13_ ( .D(n570), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[13]) );
  DFFRX1 MulCntrl_Op2_reg_14_ ( .D(n569), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[14]) );
  DFFRX1 MulCntrl_Op2_reg_15_ ( .D(n568), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[15]) );
  DFFRX1 MulCntrl_Op1_reg_0_ ( .D(n567), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[0]) );
  DFFRX1 MulCntrl_Op1_reg_1_ ( .D(n566), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[1]) );
  DFFRX1 MulCntrl_Op1_reg_2_ ( .D(n565), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[2]) );
  DFFRX1 MulCntrl_Op1_reg_3_ ( .D(n564), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[3]) );
  DFFRX1 MulCntrl_Op1_reg_4_ ( .D(n563), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[4]) );
  DFFRX1 MulCntrl_Op1_reg_5_ ( .D(n562), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[5]) );
  DFFRX1 MulCntrl_Op1_reg_6_ ( .D(n561), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[6]) );
  DFFRX1 MulCntrl_Op1_reg_7_ ( .D(n560), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[7]) );
  DFFRX1 MulCntrl_Op1_reg_8_ ( .D(n559), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[8]) );
  DFFRX1 MulCntrl_Op1_reg_9_ ( .D(n558), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[9]) );
  DFFRX1 MulCntrl_Op1_reg_10_ ( .D(n557), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[10]) );
  DFFRX1 MulCntrl_Op1_reg_11_ ( .D(n556), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[11]) );
  DFFRX1 MulCntrl_Op1_reg_12_ ( .D(n555), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[12]) );
  DFFRX1 MulCntrl_Op1_reg_13_ ( .D(n554), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[13]) );
  DFFRX1 MulCntrl_Op1_reg_14_ ( .D(n553), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[14]) );
  DFFRX1 MulCntrl_Op1_reg_15_ ( .D(n552), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[15]) );
  DFFRX1 MBUSY_reg ( .D(N150), .CLK(CLK), .CLRB(n408), .Q(MBUSY) );
  DFFRX1 DR_reg ( .D(N191), .CLK(CLK), .CLRB(n408), .Q(DR) );
  DFFRX1 MultExc_reg_reg_2_ ( .D(n469), .CLK(CLK), .CLRB(n408), .Q(
        MultExc_reg[2]) );
  DFFRX1 MultExc_reg_reg_1_ ( .D(n468), .CLK(CLK), .CLRB(n408), .Q(
        MultExc_reg[1]) );
  DFFRX1 MultExc_reg_reg_0_ ( .D(n467), .CLK(CLK), .CLRB(n408), .Q(
        MultExc_reg[0]) );
  DFFRX1 MultResult_reg_reg_0_ ( .D(n470), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[0]) );
  DFFRX1 MultResult_reg_reg_1_ ( .D(n471), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[1]) );
  DFFRX1 MultResult_reg_reg_2_ ( .D(n472), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[2]) );
  DFFRX1 MultResult_reg_reg_3_ ( .D(n473), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[3]) );
  DFFRX1 MultResult_reg_reg_4_ ( .D(n474), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[4]) );
  DFFRX1 MultResult_reg_reg_5_ ( .D(n475), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[5]) );
  DFFRX1 MultResult_reg_reg_6_ ( .D(n476), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[6]) );
  DFFRX1 MultResult_reg_reg_7_ ( .D(n477), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[7]) );
  DFFRX1 MultResult_reg_reg_8_ ( .D(n478), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[8]) );
  DFFRX1 MultResult_reg_reg_9_ ( .D(n479), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[9]) );
  DFFRX1 MultResult_reg_reg_10_ ( .D(n480), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[10]) );
  DFFRX1 MultResult_reg_reg_11_ ( .D(n481), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[11]) );
  DFFRX1 MultResult_reg_reg_12_ ( .D(n482), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[12]) );
  DFFRX1 MultResult_reg_reg_13_ ( .D(n483), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[13]) );
  DFFRX1 MultResult_reg_reg_14_ ( .D(n484), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[14]) );
  DFFRX1 MultResult_reg_reg_15_ ( .D(n485), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[15]) );
  DFFRX1 u_booth_Adder_datain1_reg_6_ ( .D(u_booth_N55), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[6]) );
  DFFRX1 u_booth_Adder_datain1_reg_7_ ( .D(n709), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain1[7]) );
  DFFRX1 u_booth_Adder_datain1_reg_8_ ( .D(n710), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain1[8]) );
  DFFRX1 u_Adder_interconnect_Select_reg ( .D(n1723), .CLK(CLK), .CLRB(n408), 
        .Q(AddSelect), .QB(n1804) );
  NANDX2 add_x_173_U10 ( .IN1(add_x_173_n64), .IN2(add_x_173_n35), .OUT(
        add_x_173_n23) );
  NANDX2 add_x_173_U77 ( .IN1(add_x_173_n71), .IN2(add_x_173_n1), .OUT(
        add_x_173_n30) );
  NANDX2 add_x_173_U13 ( .IN1(Add_Op2_wire[8]), .IN2(Add_Op1_wire[8]), .OUT(
        add_x_173_n35) );
  NANDX2 add_x_173_U26 ( .IN1(Add_Op2_wire[6]), .IN2(Add_Op1_wire[6]), .OUT(
        add_x_173_n41) );
  NANDX2 add_x_173_U35 ( .IN1(Add_Op2_wire[5]), .IN2(Add_Op1_wire[5]), .OUT(
        add_x_173_n44) );
  NANDX2 add_x_173_U66 ( .IN1(Add_Op2_wire[2]), .IN2(Add_Op1_wire[2]), .OUT(
        add_x_173_n57) );
  NANDX2 add_x_173_U55 ( .IN1(Add_Op2_wire[3]), .IN2(Add_Op1_wire[3]), .OUT(
        add_x_173_n52) );
  NANDX2 add_x_173_U75 ( .IN1(Add_Op2_wire[1]), .IN2(Add_Op1_wire[1]), .OUT(
        add_x_173_n60) );
  NANDX2 add_x_173_U80 ( .IN1(Add_Op1_wire[0]), .IN2(Add_Op2_wire[0]), .OUT(
        add_x_173_n1) );
  NANDX2 add_x_173_U46 ( .IN1(Add_Op2_wire[4]), .IN2(Add_Op1_wire[4]), .OUT(
        add_x_173_n49) );
  NOR2X1 add_x_173_U79 ( .IN1(Add_Op2_wire[0]), .IN2(Add_Op1_wire[0]), .OUT(
        add_x_173_n61) );
  NOR2X1 add_x_173_U74 ( .IN1(Add_Op1_wire[1]), .IN2(Add_Op2_wire[1]), .OUT(
        add_x_173_n59) );
  OAI21 add_x_173_U71 ( .IN1(add_x_173_n1), .IN2(add_x_173_n59), .IN3(
        add_x_173_n60), .OUT(add_x_173_n58) );
  NOR2X1 add_x_173_U65 ( .IN1(Add_Op1_wire[2]), .IN2(Add_Op2_wire[2]), .OUT(
        add_x_173_n56) );
  NOR2X1 add_x_173_U54 ( .IN1(Add_Op1_wire[3]), .IN2(Add_Op2_wire[3]), .OUT(
        add_x_173_n51) );
  NOR2X1 add_x_173_U45 ( .IN1(Add_Op1_wire[4]), .IN2(Add_Op2_wire[4]), .OUT(
        add_x_173_n48) );
  NOR2X1 add_x_173_U34 ( .IN1(Add_Op1_wire[5]), .IN2(Add_Op2_wire[5]), .OUT(
        add_x_173_n43) );
  NOR2X1 add_x_173_U25 ( .IN1(Add_Op1_wire[6]), .IN2(Add_Op2_wire[6]), .OUT(
        add_x_173_n40) );
  AOI21 add_x_173_U20 ( .IN1(add_x_173_n42), .IN2(add_x_173_n65), .IN3(
        add_x_173_n39), .OUT(add_x_173_n37) );
  FULLADD add_x_173_U14 ( .A(Add_Op2_wire[7]), .B(Add_Op1_wire[7]), .CIN(
        add_x_173_n63), .COUT(add_x_173_n36), .SUM(u_adder_24b_N129) );
  NOR2X1 add_x_173_U12 ( .IN1(Add_Op1_wire[8]), .IN2(Add_Op2_wire[8]), .OUT(
        add_x_173_n34) );
  AOI21 add_x_173_U7 ( .IN1(add_x_173_n36), .IN2(add_x_173_n64), .IN3(
        add_x_173_n33), .OUT(add_x_173_n31) );
  INVX1 U1588 ( .IN(n1802), .OUT(n1725) );
  OAI21 U1589 ( .IN1(n1801), .IN2(n1795), .IN3(n1725), .OUT(add_x_173_n42) );
  INVX1 U1590 ( .IN(add_x_173_n1), .OUT(n1726) );
  INVX1 U1591 ( .IN(add_x_173_n60), .OUT(n1727) );
  NOR2X1 U1592 ( .IN1(add_x_173_n59), .IN2(n1727), .OUT(n1728) );
  MUX2X1 U1593 ( .IN1(n1726), .IN2(add_x_173_n1), .S(n1728), .OUT(n1729) );
  AOI22 U1594 ( .IN1(Add_dataout[1]), .IN2(n2008), .IN3(n2030), .IN4(n1729), 
        .OUT(n1730) );
  INVX1 U1595 ( .IN(n1730), .OUT(n605) );
  NAND3X1 U1596 ( .IN1(add_x_173_n52), .IN2(n1797), .IN3(add_x_173_n49), .OUT(
        n1731) );
  INVX1 U1597 ( .IN(n1731), .OUT(n1798) );
  INVX1 U1598 ( .IN(add_x_173_n58), .OUT(n1732) );
  NAND2X1 U1599 ( .IN1(add_x_173_n57), .IN2(add_x_173_n69), .OUT(n1733) );
  MUX2X1 U1600 ( .IN1(n1732), .IN2(add_x_173_n58), .S(n1733), .OUT(n1734) );
  AOI22 U1601 ( .IN1(n2030), .IN2(n1734), .IN3(n2008), .IN4(Add_dataout[2]), 
        .OUT(n1735) );
  INVX1 U1602 ( .IN(n1735), .OUT(n604) );
  AOI22 U1603 ( .IN1(n2021), .IN2(n1812), .IN3(n2024), .IN4(n1841), .OUT(n1736) );
  AOI21 U1604 ( .IN1(n2022), .IN2(Add_dataout[1]), .IN3(u_booth_N49), .OUT(
        n1737) );
  NAND2X1 U1605 ( .IN1(n1736), .IN2(n1737), .OUT(n1553) );
  NAND2X1 U1606 ( .IN1(add_x_173_n52), .IN2(n1793), .OUT(n1738) );
  INVX1 U1607 ( .IN(n1738), .OUT(n1739) );
  AOI21 U1608 ( .IN1(add_x_173_n58), .IN2(add_x_173_n69), .IN3(add_x_173_n55), 
        .OUT(n1740) );
  MUX2X1 U1609 ( .IN1(n1738), .IN2(n1739), .S(n1740), .OUT(n1741) );
  AOI22 U1610 ( .IN1(Add_dataout[3]), .IN2(n2008), .IN3(n2030), .IN4(n1741), 
        .OUT(n1742) );
  INVX1 U1611 ( .IN(n1742), .OUT(n603) );
  AOI22 U1612 ( .IN1(n2021), .IN2(n1839), .IN3(n1812), .IN4(n2024), .OUT(n1743) );
  AOI21 U1613 ( .IN1(n2022), .IN2(Add_dataout[2]), .IN3(u_booth_N50), .OUT(
        n1744) );
  NAND2X1 U1614 ( .IN1(n1743), .IN2(n1744), .OUT(n1552) );
  NOR2X1 U1615 ( .IN1(add_x_173_n48), .IN2(n1745), .OUT(n1746) );
  INVX1 U1616 ( .IN(n1746), .OUT(n1747) );
  NAND3X1 U1617 ( .IN1(n1795), .IN2(n1797), .IN3(add_x_173_n52), .OUT(n1748)
         );
  MUX2X1 U1618 ( .IN1(n1746), .IN2(n1747), .S(n1748), .OUT(n1749) );
  AOI22 U1619 ( .IN1(n2030), .IN2(n1749), .IN3(n2008), .IN4(Add_dataout[4]), 
        .OUT(n1750) );
  INVX1 U1620 ( .IN(n1750), .OUT(n602) );
  INVX1 U1621 ( .IN(add_x_173_n49), .OUT(n1745) );
  AOI22 U1622 ( .IN1(n2021), .IN2(n1811), .IN3(n1839), .IN4(n2024), .OUT(n1751) );
  AOI21 U1623 ( .IN1(n2022), .IN2(Add_dataout[3]), .IN3(u_booth_N51), .OUT(
        n1752) );
  NAND2X1 U1624 ( .IN1(n1751), .IN2(n1752), .OUT(n1551) );
  NAND2X1 U1625 ( .IN1(add_x_173_n44), .IN2(n1800), .OUT(n1753) );
  INVX1 U1626 ( .IN(n1753), .OUT(n1754) );
  INVX1 U1627 ( .IN(n1796), .OUT(n1755) );
  AOI21 U1628 ( .IN1(n1795), .IN2(n1798), .IN3(n1755), .OUT(n1756) );
  MUX2X1 U1629 ( .IN1(n1754), .IN2(n1753), .S(n1756), .OUT(n1757) );
  AOI22 U1630 ( .IN1(Add_dataout[5]), .IN2(n2008), .IN3(n2030), .IN4(n1757), 
        .OUT(n1758) );
  INVX1 U1631 ( .IN(n1758), .OUT(n601) );
  NAND3X1 U1632 ( .IN1(MulCntrl_ExcCheck_Datain[10]), .IN2(ExcSelect), .IN3(
        MulCntrl_ExcCheck_Datain[7]), .OUT(n1759) );
  INVX1 U1633 ( .IN(n1759), .OUT(n1760) );
  NAND3X1 U1634 ( .IN1(MulCntrl_ExcCheck_Datain[11]), .IN2(
        MulCntrl_ExcCheck_Datain[12]), .IN3(MulCntrl_ExcCheck_Datain[13]), 
        .OUT(n1761) );
  NAND3X1 U1635 ( .IN1(MulCntrl_ExcCheck_Datain[8]), .IN2(
        MulCntrl_ExcCheck_Datain[9]), .IN3(MulCntrl_ExcCheck_Datain[14]), 
        .OUT(n1762) );
  NOR2X1 U1636 ( .IN1(n1761), .IN2(n1762), .OUT(n1763) );
  NAND3X1 U1637 ( .IN1(AdderCntrl_ExcCheck_Datain[12]), .IN2(
        AdderCntrl_ExcCheck_Datain[14]), .IN3(AdderCntrl_ExcCheck_Datain[11]), 
        .OUT(n1764) );
  NOR2X1 U1638 ( .IN1(AdderCntrl_ExcCheck_Datain[7]), .IN2(n1764), .OUT(n1765)
         );
  NOR2X1 U1639 ( .IN1(AdderCntrl_ExcCheck_Datain[13]), .IN2(
        AdderCntrl_ExcCheck_Datain[10]), .OUT(n1766) );
  NAND3X1 U1640 ( .IN1(AdderCntrl_ExcCheck_Datain[8]), .IN2(
        AdderCntrl_ExcCheck_Datain[9]), .IN3(n1766), .OUT(n1767) );
  NOR2X1 U1641 ( .IN1(ExcSelect), .IN2(n1767), .OUT(n1768) );
  AOI22 U1642 ( .IN1(n1760), .IN2(n1763), .IN3(n1765), .IN4(n1768), .OUT(n2199) );
  AOI22 U1643 ( .IN1(n2021), .IN2(n1842), .IN3(n1811), .IN4(n2024), .OUT(n1769) );
  AOI21 U1644 ( .IN1(n2022), .IN2(Add_dataout[4]), .IN3(u_booth_N52), .OUT(
        n1770) );
  NAND2X1 U1645 ( .IN1(n1769), .IN2(n1770), .OUT(n1550) );
  INVX1 U1646 ( .IN(add_x_173_n42), .OUT(n1771) );
  NAND2X1 U1647 ( .IN1(add_x_173_n41), .IN2(add_x_173_n65), .OUT(n1772) );
  MUX2X1 U1648 ( .IN1(n1771), .IN2(add_x_173_n42), .S(n1772), .OUT(n1773) );
  AOI22 U1649 ( .IN1(n2030), .IN2(n1773), .IN3(n2008), .IN4(Add_dataout[6]), 
        .OUT(n1774) );
  INVX1 U1650 ( .IN(n1774), .OUT(n600) );
  NAND3X1 U1651 ( .IN1(n714), .IN2(n1918), .IN3(u_booth_Q1_reg), .OUT(n1945)
         );
  NAND3X1 U1652 ( .IN1(u_Adder_interconnect_stateMC_1_), .IN2(n1843), .IN3(
        n806), .OUT(n1897) );
  AOI22 U1653 ( .IN1(n2026), .IN2(DIN1[13]), .IN3(MulCntrl_Op1[13]), .IN4(
        n2027), .OUT(n1775) );
  INVX1 U1654 ( .IN(n1775), .OUT(n554) );
  AOI22 U1655 ( .IN1(n2021), .IN2(n1810), .IN3(n2024), .IN4(n1842), .OUT(n1776) );
  AOI21 U1656 ( .IN1(n2022), .IN2(Add_dataout[5]), .IN3(u_booth_N53), .OUT(
        n1777) );
  NAND2X1 U1657 ( .IN1(n1776), .IN2(n1777), .OUT(n1549) );
  AOI21 U1658 ( .IN1(add_x_173_n23), .IN2(add_x_173_n36), .IN3(n1792), .OUT(
        n1778) );
  INVX1 U1659 ( .IN(n2030), .OUT(n1779) );
  NAND2X1 U1660 ( .IN1(n2008), .IN2(Add_dataout[8]), .OUT(n1780) );
  OAI21 U1661 ( .IN1(n1778), .IN2(n1779), .IN3(n1780), .OUT(n598) );
  INVX4 U1662 ( .IN(AdderCntrl_ExcCheck_Datain[7]), .OUT(n1781) );
  INVX4 U1663 ( .IN(AdderCntrl_ExcCheck_Datain[10]), .OUT(n1782) );
  INVX4 U1664 ( .IN(Booth_ack), .OUT(n1783) );
  BUF4X U1665 ( .IN(n1852), .OUT(n1784) );
  BUF4X U1666 ( .IN(AdderCntrl_Op2[8]), .OUT(n1870) );
  NAND2X1 U1667 ( .IN1(n1791), .IN2(n694), .OUT(n1785) );
  BUF4X U1668 ( .IN(n1855), .OUT(n1786) );
  INVX4 U1669 ( .IN(n1878), .OUT(n1877) );
  INVX1 U1670 ( .IN(n1854), .OUT(Booth_ack) );
  NANDX2 U1671 ( .IN1(n1791), .IN2(n694), .OUT(n1853) );
  INVX4 U1672 ( .IN(n1790), .OUT(n1791) );
  BUF8X U1673 ( .IN(Booth_dataout[8]), .OUT(n1867) );
  BUF8X U1674 ( .IN(Booth_dataout[11]), .OUT(n1866) );
  BUF4X U1675 ( .IN(n1856), .OUT(n1787) );
  NAND2X1 U1676 ( .IN1(n1951), .IN2(n1906), .OUT(n2024) );
  NAND2X1 U1677 ( .IN1(RSTn), .IN2(n1845), .OUT(n1888) );
  INVX1 U1678 ( .IN(n2203), .OUT(n588) );
  INVX1 U1679 ( .IN(n1921), .OUT(n704) );
  INVX1 U1680 ( .IN(n1924), .OUT(n703) );
  INVX1 U1681 ( .IN(n1949), .OUT(n596) );
  INVX1 U1682 ( .IN(n1933), .OUT(n699) );
  INVX1 U1683 ( .IN(n1928), .OUT(n701) );
  INVX1 U1684 ( .IN(n1930), .OUT(n700) );
  INVX1 U1685 ( .IN(n1926), .OUT(n702) );
  INVX1 U1686 ( .IN(n2254), .OUT(n480) );
  INVX1 U1687 ( .IN(n2264), .OUT(n470) );
  INVX1 U1688 ( .IN(n2233), .OUT(n537) );
  INVX1 U1689 ( .IN(n2237), .OUT(n533) );
  INVX1 U1690 ( .IN(n2239), .OUT(n531) );
  INVX1 U1691 ( .IN(n2231), .OUT(n539) );
  INVX1 U1692 ( .IN(n2236), .OUT(n534) );
  INVX1 U1693 ( .IN(n2229), .OUT(n541) );
  INVX1 U1694 ( .IN(n2252), .OUT(n482) );
  INVX1 U1695 ( .IN(n2232), .OUT(n538) );
  INVX1 U1696 ( .IN(n2255), .OUT(n479) );
  INVX1 U1697 ( .IN(n2238), .OUT(n532) );
  INVX1 U1698 ( .IN(n2230), .OUT(n540) );
  INVX1 U1699 ( .IN(n2235), .OUT(n535) );
  INVX1 U1700 ( .IN(n2234), .OUT(n536) );
  INVX1 U1701 ( .IN(n2240), .OUT(n530) );
  INVX1 U1702 ( .IN(n2262), .OUT(n472) );
  INVX1 U1703 ( .IN(n2257), .OUT(n477) );
  INVX1 U1704 ( .IN(n2253), .OUT(n481) );
  INVX1 U1705 ( .IN(n2015), .OUT(n542) );
  INVX1 U1706 ( .IN(n2241), .OUT(n529) );
  INVX1 U1707 ( .IN(n2014), .OUT(n543) );
  INVX1 U1708 ( .IN(n2016), .OUT(n528) );
  INVX1 U1709 ( .IN(n2251), .OUT(n483) );
  INVX1 U1710 ( .IN(n2017), .OUT(n527) );
  INVX1 U1711 ( .IN(n2013), .OUT(n544) );
  INVX1 U1712 ( .IN(n2256), .OUT(n478) );
  INVX1 U1713 ( .IN(n2018), .OUT(n526) );
  INVX1 U1714 ( .IN(n2228), .OUT(n545) );
  INVX1 U1715 ( .IN(n2242), .OUT(n525) );
  INVX1 U1716 ( .IN(n2261), .OUT(n473) );
  INVX1 U1717 ( .IN(n2227), .OUT(n546) );
  INVX1 U1718 ( .IN(n2226), .OUT(n547) );
  INVX1 U1719 ( .IN(n2243), .OUT(n524) );
  INVX1 U1720 ( .IN(n2225), .OUT(n548) );
  INVX1 U1721 ( .IN(n2224), .OUT(n549) );
  INVX1 U1722 ( .IN(n2260), .OUT(n474) );
  INVX1 U1723 ( .IN(n2250), .OUT(n484) );
  INVX1 U1724 ( .IN(n2223), .OUT(n550) );
  INVX1 U1725 ( .IN(n2244), .OUT(n523) );
  INVX1 U1726 ( .IN(n2222), .OUT(n551) );
  INVX1 U1727 ( .IN(n2245), .OUT(n522) );
  INVX1 U1728 ( .IN(n2249), .OUT(n485) );
  INVX1 U1729 ( .IN(n2259), .OUT(n475) );
  INVX1 U1730 ( .IN(n2246), .OUT(n521) );
  INVX1 U1731 ( .IN(n2247), .OUT(n520) );
  INVX1 U1732 ( .IN(n2258), .OUT(n476) );
  INVX1 U1733 ( .IN(n2263), .OUT(n471) );
  INVX1 U1734 ( .IN(n2209), .OUT(n579) );
  INVX1 U1735 ( .IN(n2005), .OUT(n555) );
  INVX1 U1736 ( .IN(n1996), .OUT(n572) );
  INVX1 U1737 ( .IN(n1997), .OUT(n571) );
  INVX1 U1738 ( .IN(n2004), .OUT(n556) );
  INVX1 U1739 ( .IN(n2208), .OUT(n580) );
  INVX1 U1740 ( .IN(n2207), .OUT(n581) );
  INVX1 U1741 ( .IN(n2003), .OUT(n557) );
  NAND2X1 U1742 ( .IN1(n1978), .IN2(n1975), .OUT(n1977) );
  INVX1 U1743 ( .IN(n1998), .OUT(n570) );
  INVX1 U1744 ( .IN(n2206), .OUT(n582) );
  INVX1 U1745 ( .IN(n2002), .OUT(n558) );
  INVX1 U1746 ( .IN(n1992), .OUT(n576) );
  INVX1 U1747 ( .IN(n2205), .OUT(n583) );
  INVX1 U1748 ( .IN(n2001), .OUT(n559) );
  INVX1 U1749 ( .IN(n1999), .OUT(n569) );
  INVX1 U1750 ( .IN(n2000), .OUT(n560) );
  INVX1 U1751 ( .IN(n2219), .OUT(n561) );
  INVX1 U1752 ( .IN(n2212), .OUT(n568) );
  INVX1 U1753 ( .IN(n2218), .OUT(n562) );
  NAND2X1 U1754 ( .IN1(n2029), .IN2(n2152), .OUT(n1546) );
  INVX1 U1755 ( .IN(n2217), .OUT(n563) );
  INVX1 U1756 ( .IN(n2213), .OUT(n567) );
  INVX1 U1757 ( .IN(n2216), .OUT(n564) );
  INVX1 U1758 ( .IN(n2215), .OUT(n565) );
  INVX1 U1759 ( .IN(n2214), .OUT(n566) );
  INVX1 U1760 ( .IN(n2211), .OUT(n577) );
  INVX1 U1761 ( .IN(n1994), .OUT(n574) );
  INVX1 U1762 ( .IN(n2269), .OUT(n467) );
  INVX1 U1763 ( .IN(n2266), .OUT(n468) );
  INVX1 U1764 ( .IN(n2210), .OUT(n578) );
  INVX1 U1765 ( .IN(n1993), .OUT(n575) );
  INVX1 U1766 ( .IN(n2265), .OUT(n469) );
  INVX1 U1767 ( .IN(n1995), .OUT(n573) );
  INVX1 U1768 ( .IN(n2220), .OUT(n552) );
  INVX1 U1769 ( .IN(n2006), .OUT(n553) );
  NANDX2 U1770 ( .IN1(n1810), .IN2(n2023), .OUT(n2148) );
  NANDX2 U1771 ( .IN1(n1851), .IN2(n2023), .OUT(n2150) );
  INVX1 U1772 ( .IN(n2286), .OUT(n416) );
  INVX1 U1773 ( .IN(n2272), .OUT(n430) );
  INVX1 U1774 ( .IN(n2273), .OUT(n429) );
  INVX1 U1775 ( .IN(n2274), .OUT(n428) );
  NAND2X1 U1776 ( .IN1(n2113), .IN2(n2112), .OUT(n2114) );
  INVX1 U1777 ( .IN(n2275), .OUT(n427) );
  INVX1 U1778 ( .IN(n2276), .OUT(n426) );
  INVX1 U1779 ( .IN(n2277), .OUT(n425) );
  INVX1 U1780 ( .IN(n2278), .OUT(n424) );
  INVX1 U1781 ( .IN(n2279), .OUT(n423) );
  INVX1 U1782 ( .IN(n2280), .OUT(n422) );
  INVX1 U1783 ( .IN(n2281), .OUT(n421) );
  INVX1 U1784 ( .IN(n2288), .OUT(n414) );
  INVX1 U1785 ( .IN(n2282), .OUT(n420) );
  INVX1 U1786 ( .IN(n2289), .OUT(n413) );
  INVX1 U1787 ( .IN(n2283), .OUT(n419) );
  INVX1 U1788 ( .IN(n2292), .OUT(n412) );
  INVX1 U1789 ( .IN(n2284), .OUT(n418) );
  INVX1 U1790 ( .IN(n2287), .OUT(n415) );
  INVX1 U1791 ( .IN(n2285), .OUT(n417) );
  BUF4X U1792 ( .IN(Booth_dataout[6]), .OUT(n1868) );
  INVX1 U1793 ( .IN(add_x_173_n41), .OUT(add_x_173_n39) );
  NAND2X1 U1794 ( .IN1(n2020), .IN2(n2019), .OUT(n2023) );
  INVX1 U1795 ( .IN(add_x_173_n61), .OUT(add_x_173_n71) );
  INVX1 U1796 ( .IN(add_x_173_n35), .OUT(add_x_173_n33) );
  INVX1 U1797 ( .IN(n2181), .OUT(n615) );
  INVX1 U1798 ( .IN(n1939), .OUT(n610) );
  INVX1 U1799 ( .IN(n1938), .OUT(n609) );
  INVX1 U1800 ( .IN(n2147), .OUT(n1587) );
  INVX1 U1801 ( .IN(n2180), .OUT(n616) );
  INVX1 U1802 ( .IN(n2024), .OUT(n2020) );
  INVX1 U1803 ( .IN(n2184), .OUT(n612) );
  INVX1 U1804 ( .IN(n2183), .OUT(n613) );
  NANDX2 U1805 ( .IN1(n1808), .IN2(n1914), .OUT(n1915) );
  INVX1 U1806 ( .IN(n2185), .OUT(n611) );
  INVX1 U1807 ( .IN(n2182), .OUT(n614) );
  INVX1 U1808 ( .IN(n2031), .OUT(DEBUG[4]) );
  INVX1 U1809 ( .IN(n2033), .OUT(DEBUG[2]) );
  INVX1 U1810 ( .IN(n2041), .OUT(DEBUG[0]) );
  INVX1 U1811 ( .IN(n2046), .OUT(DEBUG[1]) );
  INVX1 U1812 ( .IN(n2051), .OUT(DOUT[13]) );
  INVX1 U1813 ( .IN(n2064), .OUT(EXC[0]) );
  INVX1 U1814 ( .IN(n2039), .OUT(DACK) );
  INVX1 U1815 ( .IN(n2050), .OUT(DOUT[12]) );
  INVX1 U1816 ( .IN(n2087), .OUT(n2088) );
  INVX1 U1817 ( .IN(n2052), .OUT(DOUT[14]) );
  INVX1 U1818 ( .IN(n2053), .OUT(DOUT[15]) );
  INVX1 U1819 ( .IN(n2065), .OUT(EXC[1]) );
  INVX1 U1820 ( .IN(n2058), .OUT(DOUT[5]) );
  INVX1 U1821 ( .IN(n2059), .OUT(DOUT[6]) );
  INVX1 U1822 ( .IN(n2060), .OUT(DOUT[7]) );
  INVX1 U1823 ( .IN(n2057), .OUT(DOUT[4]) );
  INVX1 U1824 ( .IN(n2056), .OUT(DOUT[3]) );
  INVX1 U1825 ( .IN(n2055), .OUT(DOUT[2]) );
  INVX1 U1826 ( .IN(n2061), .OUT(DOUT[8]) );
  INVX1 U1827 ( .IN(n2054), .OUT(DOUT[1]) );
  INVX1 U1828 ( .IN(n2047), .OUT(DOUT[0]) );
  INVX1 U1829 ( .IN(n2062), .OUT(DOUT[9]) );
  INVX1 U1830 ( .IN(n2048), .OUT(DOUT[10]) );
  INVX1 U1831 ( .IN(n2063), .OUT(DOV) );
  INVX1 U1832 ( .IN(n2067), .OUT(EXC[2]) );
  INVX1 U1833 ( .IN(n2049), .OUT(DOUT[11]) );
  NAND2X1 U1834 ( .IN1(n2043), .IN2(AdderCntrl_Debug[2]), .OUT(n2033) );
  INVX1 U1835 ( .IN(n2032), .OUT(DEBUG[3]) );
  NAND2X1 U1836 ( .IN1(n2043), .IN2(AdderCntrl_Debug[4]), .OUT(n2031) );
  NAND2X1 U1837 ( .IN1(n1787), .IN2(n1895), .OUT(n1882) );
  INVX1 U1838 ( .IN(n1887), .OUT(n1588) );
  INVX1 U1839 ( .IN(n2105), .OUT(n1656) );
  INVX1 U1840 ( .IN(n2191), .OUT(n594) );
  NANDX2 U1841 ( .IN1(Booth_Add_datain1[8]), .IN2(n1946), .OUT(n1899) );
  INVX1 U1842 ( .IN(n2196), .OUT(n592) );
  NAND2X1 U1843 ( .IN1(n2043), .IN2(AdderCntrl_Debug[3]), .OUT(n2032) );
  INVX1 U1844 ( .IN(n1904), .OUT(n1905) );
  INVX1 U1845 ( .IN(n1892), .OUT(n1893) );
  INVX1 U1846 ( .IN(n1859), .OUT(n1858) );
  INVX1 U1847 ( .IN(n2200), .OUT(n2201) );
  NANDX2 U1848 ( .IN1(Add_Op2[7]), .IN2(n1947), .OUT(n1922) );
  NAND2X1 U1849 ( .IN1(n2076), .IN2(n2086), .OUT(n2077) );
  NANDX2 U1850 ( .IN1(n1808), .IN2(n1895), .OUT(n1953) );
  INVX1 U1851 ( .IN(n2192), .OUT(n2194) );
  INVX1 U1852 ( .IN(n1888), .OUT(n1885) );
  INVX1 U1853 ( .IN(n2187), .OUT(n2190) );
  INVX1 U1854 ( .IN(n2161), .OUT(n2104) );
  NAND2X1 U1855 ( .IN1(RSTn), .IN2(n1935), .OUT(n1936) );
  NAND2X1 U1856 ( .IN1(n1860), .IN2(n1819), .OUT(n1859) );
  NANDX2 U1857 ( .IN1(multStateMC[0]), .IN2(n1807), .OUT(n2156) );
  NANDX2 U1858 ( .IN1(n1878), .IN2(n768), .OUT(n1879) );
  BUF4X U1859 ( .IN(AdderCntrl_Op1[9]), .OUT(n1869) );
  INVX4 U1860 ( .IN(CS), .OUT(n2086) );
  INVX1 U1861 ( .IN(n1788), .OUT(n1789) );
  NOR2X1 U1862 ( .IN1(add_x_173_n23), .IN2(add_x_173_n36), .OUT(n1792) );
  OAI21 U1863 ( .IN1(n1801), .IN2(n1798), .IN3(add_x_173_n44), .OUT(n1802) );
  INVX1 U1864 ( .IN(add_x_173_n43), .OUT(n1800) );
  INVX1 U1865 ( .IN(add_x_173_n40), .OUT(add_x_173_n65) );
  NANDX2 U1866 ( .IN1(add_x_173_n49), .IN2(add_x_173_n48), .OUT(n1796) );
  INVX4 U1867 ( .IN(add_x_173_n57), .OUT(add_x_173_n55) );
  NANDX2 U1868 ( .IN1(add_x_173_n55), .IN2(n1793), .OUT(n1797) );
  INVX4 U1869 ( .IN(add_x_173_n37), .OUT(add_x_173_n63) );
  INVX4 U1870 ( .IN(add_x_173_n30), .OUT(u_adder_24b_N122) );
  INVX4 U1871 ( .IN(add_x_173_n51), .OUT(n1793) );
  NANDX2 U1872 ( .IN1(add_x_173_n58), .IN2(n1799), .OUT(n1795) );
  INVX4 U1873 ( .IN(add_x_173_n56), .OUT(add_x_173_n69) );
  NANDX2 U1874 ( .IN1(n1793), .IN2(add_x_173_n69), .OUT(n1794) );
  INVX4 U1875 ( .IN(n1794), .OUT(n1799) );
  NANDX2 U1876 ( .IN1(n1800), .IN2(n1796), .OUT(n1801) );
  INVX4 U1877 ( .IN(add_x_173_n34), .OUT(add_x_173_n64) );
  INVX1 U1878 ( .IN(add_x_173_n31), .OUT(u_adder_24b_N131) );
  BUF8X U1879 ( .IN(Booth_dataout[10]), .OUT(n1864) );
  BUF4X U1880 ( .IN(n1855), .OUT(n1854) );
  INVX4 U1881 ( .IN(n1953), .OUT(n1883) );
  INVX4 U1882 ( .IN(n1952), .OUT(n1970) );
  NAND2X1 U1883 ( .IN1(n2108), .IN2(n2107), .OUT(n2109) );
  INVX4 U1884 ( .IN(n1991), .OUT(n2026) );
  INVX4 U1885 ( .IN(n2012), .OUT(n1876) );
  NANDX2 U1886 ( .IN1(n1878), .IN2(n2159), .OUT(n992) );
  NANDX2 U1887 ( .IN1(n2151), .IN2(n2150), .OUT(n1547) );
  NANDX2 U1888 ( .IN1(n2149), .IN2(n2148), .OUT(n1548) );
  INVX4 U1889 ( .IN(n2011), .OUT(n2025) );
  BUF4X U1890 ( .IN(n2267), .OUT(n1874) );
  BUF4X U1891 ( .IN(n2290), .OUT(n1875) );
  INVX4 U1892 ( .IN(n1923), .OUT(n1946) );
  INVX4 U1893 ( .IN(n1897), .OUT(n2146) );
  INVX4 U1894 ( .IN(n1990), .OUT(n2027) );
  INVX4 U1895 ( .IN(n2082), .OUT(n2268) );
  BUF4X U1896 ( .IN(n2066), .OUT(n1873) );
  NANDX2 U1897 ( .IN1(n1878), .IN2(n2090), .OUT(n1302) );
  BUF4X U1898 ( .IN(n2080), .OUT(n1872) );
  INVX4 U1899 ( .IN(n2270), .OUT(n2291) );
  NANDX2 U1900 ( .IN1(u_exc_check_N45), .IN2(n2133), .OUT(n2134) );
  NANDX2 U1901 ( .IN1(n1878), .IN2(n2106), .OUT(n2200) );
  NAND2X1 U1902 ( .IN1(n1878), .IN2(n1843), .OUT(n2137) );
  NAND2X1 U1903 ( .IN1(n1878), .IN2(u_booth_BStateMC_1_), .OUT(n1951) );
  NANDX2 U1904 ( .IN1(n1813), .IN2(n1900), .OUT(n1923) );
  NAND2X1 U1905 ( .IN1(u_booth_M_reg_1_), .IN2(n1940), .OUT(n1941) );
  INVX4 U1906 ( .IN(n1954), .OUT(n1969) );
  NANDX2 U1907 ( .IN1(n1878), .IN2(n1990), .OUT(n1991) );
  NANDX2 U1908 ( .IN1(n1878), .IN2(n1989), .OUT(n1990) );
  NAND2X1 U1909 ( .IN1(n734), .IN2(n1937), .OUT(n1952) );
  INVX1 U1910 ( .IN(Booth_valid), .OUT(n2135) );
  NANDX2 U1911 ( .IN1(RSTn), .IN2(n2011), .OUT(n2012) );
  NANDX2 U1912 ( .IN1(n1878), .IN2(n2010), .OUT(n2011) );
  NANDX2 U1913 ( .IN1(n1914), .IN2(n1893), .OUT(n1894) );
  NAND2X1 U1914 ( .IN1(n587), .IN2(CS), .OUT(n2078) );
  NAND2X1 U1915 ( .IN1(CS), .IN2(n2268), .OUT(n2155) );
  NANDX2 U1916 ( .IN1(n1878), .IN2(n2248), .OUT(n2082) );
  INVX4 U1917 ( .IN(MulCntrl_Dataout_valid), .OUT(n2079) );
  NANDX2 U1918 ( .IN1(n1878), .IN2(n2271), .OUT(n2270) );
  NANDX2 U1919 ( .IN1(n1913), .IN2(n1912), .OUT(n1984) );
  NANDX2 U1920 ( .IN1(n1914), .IN2(n1896), .OUT(n1912) );
  NAND2X1 U1921 ( .IN1(n1846), .IN2(n1914), .OUT(n1913) );
  INVX4 U1922 ( .IN(n1983), .OUT(n1975) );
  INVX4 U1923 ( .IN(n1882), .OUT(n1890) );
  NANDX2 U1924 ( .IN1(n1916), .IN2(n1918), .OUT(n1944) );
  INVX4 U1925 ( .IN(n1915), .OUT(n1918) );
  NANDX2 U1926 ( .IN1(n1878), .IN2(n1787), .OUT(n1988) );
  INVX4 U1927 ( .IN(n2198), .OUT(n2132) );
  NANDX2 U1928 ( .IN1(n2122), .IN2(n2127), .OUT(n2198) );
  INVX4 U1929 ( .IN(n1917), .OUT(Add_Op2_wire[8]) );
  INVX4 U1930 ( .IN(n1899), .OUT(Add_Op1_wire[8]) );
  INVX4 U1931 ( .IN(n1925), .OUT(Add_Op2_wire[6]) );
  INVX4 U1932 ( .IN(n1902), .OUT(Add_Op1_wire[6]) );
  INVX4 U1933 ( .IN(n1934), .OUT(Add_Op2_wire[2]) );
  INVX4 U1934 ( .IN(n1909), .OUT(Add_Op1_wire[2]) );
  INVX4 U1935 ( .IN(n1931), .OUT(Add_Op2_wire[3]) );
  INVX4 U1936 ( .IN(n1908), .OUT(Add_Op1_wire[3]) );
  INVX4 U1937 ( .IN(n1943), .OUT(Add_Op2_wire[1]) );
  INVX4 U1938 ( .IN(n1910), .OUT(Add_Op1_wire[1]) );
  INVX4 U1939 ( .IN(n1948), .OUT(Add_Op2_wire[0]) );
  INVX4 U1940 ( .IN(n1911), .OUT(Add_Op1_wire[0]) );
  INVX4 U1941 ( .IN(n1907), .OUT(Add_Op1_wire[4]) );
  INVX4 U1942 ( .IN(n1929), .OUT(Add_Op2_wire[4]) );
  INVX4 U1943 ( .IN(n1927), .OUT(Add_Op2_wire[5]) );
  INVX4 U1944 ( .IN(n1903), .OUT(Add_Op1_wire[5]) );
  INVX4 U1945 ( .IN(n1901), .OUT(Add_Op1_wire[7]) );
  INVX4 U1946 ( .IN(n1879), .OUT(n1880) );
  NANDX2 U1947 ( .IN1(n1889), .IN2(n1888), .OUT(n2008) );
  INVX4 U1948 ( .IN(n1803), .OUT(n1871) );
  INVX4 U1949 ( .IN(n1857), .OUT(Booth_dataout[12]) );
  INVX4 U1950 ( .IN(n1861), .OUT(n1852) );
  BUF4X U1951 ( .IN(RSTn), .OUT(n1878) );
  NAND2X1 U1952 ( .IN1(n1846), .IN2(n1895), .OUT(n1892) );
  NAND2X1 U1953 ( .IN1(n1878), .IN2(n1838), .OUT(n1884) );
  INVX1 U1954 ( .IN(n2176), .OUT(n2175) );
  NAND2X1 U1955 ( .IN1(n1905), .IN2(n734), .OUT(n1906) );
  NAND2X1 U1956 ( .IN1(n2135), .IN2(n1878), .OUT(n1904) );
  INVX1 U1957 ( .IN(n2204), .OUT(n1989) );
  NAND2X1 U1958 ( .IN1(Booth_valid), .IN2(n734), .OUT(n1935) );
  INVX1 U1959 ( .IN(n2221), .OUT(n2010) );
  NAND2X1 U1960 ( .IN1(u_booth_count_reg_2_), .IN2(n1983), .OUT(n1979) );
  NAND2X1 U1961 ( .IN1(u_booth_count_reg_2_), .IN2(n1978), .OUT(n1982) );
  INVX1 U1962 ( .IN(n1895), .OUT(n1896) );
  NAND2X1 U1963 ( .IN1(u_booth_M_reg_7_), .IN2(n1919), .OUT(n1920) );
  INVX1 U1964 ( .IN(n2162), .OUT(n1919) );
  INVX1 U1965 ( .IN(n2009), .OUT(n599) );
  INVX1 U1966 ( .IN(n2007), .OUT(n597) );
  NAND2X1 U1967 ( .IN1(RSTn), .IN2(u_adder_24b_StateMC_1_), .OUT(n1889) );
  BUF4X U1968 ( .IN(MulCntrl_Op2[8]), .OUT(n1862) );
  BUF4X U1969 ( .IN(MulCntrl_Op1[8]), .OUT(n1865) );
  BUF4X U1970 ( .IN(MulCntrl_Op2[13]), .OUT(n1863) );
  NAND2X1 U1971 ( .IN1(n1852), .IN2(n1858), .OUT(n1857) );
  NANDX2 U1972 ( .IN1(n1787), .IN2(n1852), .OUT(n1855) );
  OAI21 U1973 ( .IN1(n1988), .IN2(n1784), .IN3(n1987), .OUT(n1556) );
  OAI21 U1974 ( .IN1(u_booth_count_reg_2_), .IN2(n1853), .IN3(
        u_booth_count_reg_3_), .OUT(n1861) );
  NAND3X1 U1975 ( .IN1(n1977), .IN2(n1785), .IN3(n1976), .OUT(n1080) );
  NOR2X1 U1976 ( .IN1(u_booth_BStateMC_1_), .IN2(n1789), .OUT(n1856) );
  NOR2X1 U1977 ( .IN1(n722), .IN2(n1855), .OUT(Booth_dataout[8]) );
  NOR2X1 U1978 ( .IN1(n721), .IN2(n1855), .OUT(Booth_dataout[7]) );
  NOR2X1 U1979 ( .IN1(n724), .IN2(n1855), .OUT(Booth_dataout[10]) );
  NOR2X1 U1980 ( .IN1(n723), .IN2(n1855), .OUT(Booth_dataout[9]) );
  NOR2X1 U1981 ( .IN1(n720), .IN2(n1855), .OUT(Booth_dataout[6]) );
  NOR2X1 U1982 ( .IN1(n725), .IN2(n1855), .OUT(Booth_dataout[11]) );
  NOR2X1 U1983 ( .IN1(n727), .IN2(n1855), .OUT(Booth_dataout[13]) );
  NOR2X1 U1984 ( .IN1(n717), .IN2(n1855), .OUT(Booth_dataout[3]) );
  NOR2X1 U1985 ( .IN1(n714), .IN2(n1854), .OUT(Booth_dataout[0]) );
  NOR2X1 U1986 ( .IN1(n729), .IN2(n1854), .OUT(Booth_dataout[15]) );
  NOR2X1 U1987 ( .IN1(n728), .IN2(n1783), .OUT(Booth_dataout[14]) );
  NAND2X1 U1988 ( .IN1(n1787), .IN2(n1953), .OUT(n1954) );
  NOR2X1 U1989 ( .IN1(n726), .IN2(n734), .OUT(n1860) );
  TIELO U1990 ( .OUT(n2293) );
  TIEHI U1991 ( .OUT(n408) );
  NOR2X1 U1992 ( .IN1(n734), .IN2(n1951), .OUT(n1986) );
  AOI21 U1993 ( .IN1(Booth_ack), .IN2(RSTn), .IN3(n1986), .OUT(n1089) );
  NOR2X1 U1994 ( .IN1(n802), .IN2(u_adder_24b_StateMC_1_), .OUT(n1886) );
  NANDX2 U1995 ( .IN1(n1880), .IN2(n1886), .OUT(n1881) );
  INVX4 U1996 ( .IN(n1881), .OUT(n2030) );
  AOI22 U1997 ( .IN1(n1816), .IN2(n714), .IN3(u_booth_Q1_reg), .IN4(n1806), 
        .OUT(n1895) );
  INVX4 U1998 ( .IN(n1988), .OUT(n1914) );
  NANDX2 U1999 ( .IN1(n1914), .IN2(n1883), .OUT(n2019) );
  OAI21 U2000 ( .IN1(n1890), .IN2(n2137), .IN3(n2019), .OUT(n1653) );
  NAND3X1 U2001 ( .IN1(Add_valid), .IN2(n1809), .IN3(n1822), .OUT(n2187) );
  AOI21 U2002 ( .IN1(n2187), .IN2(n1897), .IN3(n1884), .OUT(
        u_Adder_interconnect_N53) );
  NOR2X1 U2003 ( .IN1(n1886), .IN2(n1888), .OUT(n1589) );
  AOI22 U2004 ( .IN1(n1886), .IN2(RSTn), .IN3(u_adder_24b_StateMC_1_), .IN4(
        n1885), .OUT(n1887) );
  NOR2X1 U2005 ( .IN1(Booth_valid), .IN2(u_booth_BStateMC_1_), .OUT(n1891) );
  AOI22 U2006 ( .IN1(n1891), .IN2(n734), .IN3(n1808), .IN4(n1890), .OUT(n1972)
         );
  AOI21 U2007 ( .IN1(n1972), .IN2(n1819), .IN3(n1877), .OUT(n1983) );
  INVX4 U2008 ( .IN(n1894), .OUT(n2022) );
  INVX4 U2009 ( .IN(n1912), .OUT(n2021) );
  AOI22 U2010 ( .IN1(n2022), .IN2(Add_dataout[8]), .IN3(n2021), .IN4(
        u_booth_A_reg_8_), .OUT(n2029) );
  OAI21 U2011 ( .IN1(n1849), .IN2(n1975), .IN3(n2029), .OUT(n1545) );
  NOR2X1 U2012 ( .IN1(n1849), .IN2(n2019), .OUT(n710) );
  AOI21 U2013 ( .IN1(n2187), .IN2(AddSelect), .IN3(n2146), .OUT(n1898) );
  NOR2X1 U2014 ( .IN1(n1877), .IN2(n1898), .OUT(n1723) );
  NANDX2 U2015 ( .IN1(n1804), .IN2(n1813), .OUT(n1900) );
  NOR2X1 U2016 ( .IN1(n1828), .IN2(n2019), .OUT(n709) );
  INVX4 U2017 ( .IN(n1900), .OUT(n1947) );
  AOI22 U2018 ( .IN1(n1947), .IN2(Add_Op1[7]), .IN3(Booth_Add_datain1[7]), 
        .IN4(n1946), .OUT(n1901) );
  NOR2X1 U2019 ( .IN1(n729), .IN2(n2019), .OUT(u_booth_N55) );
  AOI22 U2020 ( .IN1(n1947), .IN2(Add_Op1[6]), .IN3(Booth_Add_datain1[6]), 
        .IN4(n1946), .OUT(n1902) );
  NOR2X1 U2021 ( .IN1(n728), .IN2(n2019), .OUT(u_booth_N54) );
  AOI22 U2022 ( .IN1(n1947), .IN2(Add_Op1[5]), .IN3(Booth_Add_datain1[5]), 
        .IN4(n1946), .OUT(n1903) );
  NOR2X1 U2023 ( .IN1(n727), .IN2(n2019), .OUT(u_booth_N53) );
  AOI22 U2024 ( .IN1(n1947), .IN2(Add_Op1[4]), .IN3(Booth_Add_datain1[4]), 
        .IN4(n1946), .OUT(n1907) );
  NOR2X1 U2025 ( .IN1(n726), .IN2(n2019), .OUT(u_booth_N52) );
  AOI22 U2026 ( .IN1(n1947), .IN2(Add_Op1[3]), .IN3(Booth_Add_datain1[3]), 
        .IN4(n1946), .OUT(n1908) );
  NOR2X1 U2027 ( .IN1(n725), .IN2(n2019), .OUT(u_booth_N51) );
  AOI22 U2028 ( .IN1(n1947), .IN2(Add_Op1[2]), .IN3(Booth_Add_datain1[2]), 
        .IN4(n1946), .OUT(n1909) );
  NOR2X1 U2029 ( .IN1(n724), .IN2(n2019), .OUT(u_booth_N50) );
  AOI22 U2030 ( .IN1(n1947), .IN2(Add_Op1[1]), .IN3(Booth_Add_datain1[1]), 
        .IN4(n1946), .OUT(n1910) );
  NOR2X1 U2031 ( .IN1(n723), .IN2(n2019), .OUT(u_booth_N49) );
  AOI22 U2032 ( .IN1(n1947), .IN2(Add_Op1[0]), .IN3(Booth_Add_datain1[0]), 
        .IN4(n1946), .OUT(n1911) );
  AOI22 U2033 ( .IN1(n1806), .IN2(n1984), .IN3(u_booth_Q1_reg), .IN4(n1983), 
        .OUT(n1078) );
  NOR2X1 U2034 ( .IN1(u_booth_Q1_reg), .IN2(n714), .OUT(n1916) );
  AOI21 U2035 ( .IN1(n2162), .IN2(n1829), .IN3(n1944), .OUT(n705) );
  AOI22 U2036 ( .IN1(n1947), .IN2(Add_Op2[8]), .IN3(Booth_Add_datain2[8]), 
        .IN4(n1946), .OUT(n1917) );
  INVX4 U2037 ( .IN(n1945), .OUT(n1940) );
  AOI22 U2038 ( .IN1(n1940), .IN2(u_booth_M_reg_7_), .IN3(n1920), .IN4(n705), 
        .OUT(n1921) );
  OAI21 U2039 ( .IN1(n1818), .IN2(n1923), .IN3(n1922), .OUT(Add_Op2_wire[7])
         );
  INVX4 U2040 ( .IN(n1944), .OUT(n1932) );
  AOI22 U2041 ( .IN1(n1940), .IN2(u_booth_M_reg_6_), .IN3(n1932), .IN4(n2165), 
        .OUT(n1924) );
  AOI22 U2042 ( .IN1(n1947), .IN2(Add_Op2[6]), .IN3(Booth_Add_datain2[6]), 
        .IN4(n1946), .OUT(n1925) );
  AOI22 U2043 ( .IN1(n1940), .IN2(u_booth_M_reg_5_), .IN3(n1932), .IN4(n2168), 
        .OUT(n1926) );
  AOI22 U2044 ( .IN1(n1947), .IN2(Add_Op2[5]), .IN3(Booth_Add_datain2[5]), 
        .IN4(n1946), .OUT(n1927) );
  AOI22 U2045 ( .IN1(n1940), .IN2(u_booth_M_reg_4_), .IN3(n1932), .IN4(n2171), 
        .OUT(n1928) );
  AOI22 U2046 ( .IN1(n1947), .IN2(Add_Op2[4]), .IN3(Booth_Add_datain2[4]), 
        .IN4(n1946), .OUT(n1929) );
  AOI22 U2047 ( .IN1(n1940), .IN2(u_booth_M_reg_3_), .IN3(n1932), .IN4(n2174), 
        .OUT(n1930) );
  AOI22 U2048 ( .IN1(n1947), .IN2(Add_Op2[3]), .IN3(Booth_Add_datain2[3]), 
        .IN4(n1946), .OUT(n1931) );
  AOI22 U2049 ( .IN1(n1940), .IN2(u_booth_M_reg_2_), .IN3(n1932), .IN4(n2177), 
        .OUT(n1933) );
  AOI22 U2050 ( .IN1(n1947), .IN2(Add_Op2[2]), .IN3(Booth_Add_datain2[2]), 
        .IN4(n1946), .OUT(n1934) );
  NANDX2 U2051 ( .IN1(n1951), .IN2(n1936), .OUT(n2186) );
  NOR2X1 U2052 ( .IN1(n2135), .IN2(u_booth_BStateMC_1_), .OUT(n1937) );
  NOR2X1 U2053 ( .IN1(n1877), .IN2(n1952), .OUT(n2028) );
  AOI22 U2054 ( .IN1(u_booth_N258), .IN2(n2186), .IN3(Booth_datain1[0]), .IN4(
        n2028), .OUT(n1938) );
  AOI22 U2055 ( .IN1(u_booth_M_reg_1_), .IN2(n2186), .IN3(Booth_datain1[1]), 
        .IN4(n2028), .OUT(n1939) );
  AOI22 U2056 ( .IN1(n1814), .IN2(u_booth_M_reg_1_), .IN3(u_booth_N258), .IN4(
        n1805), .OUT(n1942) );
  OAI21 U2057 ( .IN1(n1942), .IN2(n1944), .IN3(n1941), .OUT(n698) );
  AOI22 U2058 ( .IN1(n1947), .IN2(Add_Op2[1]), .IN3(Booth_Add_datain2[1]), 
        .IN4(n1946), .OUT(n1943) );
  AOI21 U2059 ( .IN1(n1945), .IN2(n1944), .IN3(n1814), .OUT(n697) );
  AOI22 U2060 ( .IN1(n1947), .IN2(Add_Op2[0]), .IN3(Booth_Add_datain2[0]), 
        .IN4(n1946), .OUT(n1948) );
  AOI22 U2061 ( .IN1(Add_dataout[0]), .IN2(n2008), .IN3(n2030), .IN4(
        u_adder_24b_N122), .OUT(n1949) );
  AOI22 U2062 ( .IN1(n2021), .IN2(n1841), .IN3(Add_dataout[0]), .IN4(n2022), 
        .OUT(n1950) );
  OAI21 U2063 ( .IN1(n722), .IN2(n1975), .IN3(n1950), .OUT(n1544) );
  INVX4 U2064 ( .IN(n1951), .OUT(n1974) );
  AOI22 U2065 ( .IN1(Booth_datain2[7]), .IN2(n1970), .IN3(n1844), .IN4(n1969), 
        .OUT(n1955) );
  OAI21 U2066 ( .IN1(n721), .IN2(n1972), .IN3(n1955), .OUT(n1956) );
  AOI22 U2067 ( .IN1(n1974), .IN2(n1830), .IN3(RSTn), .IN4(n1956), .OUT(n1021)
         );
  AOI22 U2068 ( .IN1(Booth_datain2[6]), .IN2(n1970), .IN3(n1830), .IN4(n1969), 
        .OUT(n1957) );
  OAI21 U2069 ( .IN1(n720), .IN2(n1972), .IN3(n1957), .OUT(n1958) );
  AOI22 U2070 ( .IN1(n1974), .IN2(n1831), .IN3(n1878), .IN4(n1958), .OUT(n1028) );
  AOI22 U2071 ( .IN1(n1970), .IN2(Booth_datain2[5]), .IN3(n1831), .IN4(n1969), 
        .OUT(n1959) );
  OAI21 U2072 ( .IN1(n719), .IN2(n1972), .IN3(n1959), .OUT(n1960) );
  AOI22 U2073 ( .IN1(n1974), .IN2(n1832), .IN3(n1878), .IN4(n1960), .OUT(n1031) );
  AOI22 U2074 ( .IN1(n1970), .IN2(Booth_datain2[4]), .IN3(n1832), .IN4(n1969), 
        .OUT(n1961) );
  OAI21 U2075 ( .IN1(n718), .IN2(n1972), .IN3(n1961), .OUT(n1962) );
  AOI22 U2076 ( .IN1(n1974), .IN2(n1833), .IN3(n1878), .IN4(n1962), .OUT(n1034) );
  AOI22 U2077 ( .IN1(n1970), .IN2(Booth_datain2[3]), .IN3(n1833), .IN4(n1969), 
        .OUT(n1963) );
  OAI21 U2078 ( .IN1(n717), .IN2(n1972), .IN3(n1963), .OUT(n1964) );
  AOI22 U2079 ( .IN1(n1974), .IN2(n1834), .IN3(RSTn), .IN4(n1964), .OUT(n1037)
         );
  AOI22 U2080 ( .IN1(n1970), .IN2(Booth_datain2[2]), .IN3(n1834), .IN4(n1969), 
        .OUT(n1965) );
  OAI21 U2081 ( .IN1(n716), .IN2(n1972), .IN3(n1965), .OUT(n1966) );
  AOI22 U2082 ( .IN1(n1974), .IN2(n1835), .IN3(n1878), .IN4(n1966), .OUT(n1040) );
  AOI22 U2083 ( .IN1(n1970), .IN2(Booth_datain2[1]), .IN3(n1835), .IN4(n1969), 
        .OUT(n1967) );
  OAI21 U2084 ( .IN1(n715), .IN2(n1972), .IN3(n1967), .OUT(n1968) );
  AOI22 U2085 ( .IN1(n1974), .IN2(n1836), .IN3(RSTn), .IN4(n1968), .OUT(n1043)
         );
  AOI22 U2086 ( .IN1(n1970), .IN2(Booth_datain2[0]), .IN3(n1836), .IN4(n1969), 
        .OUT(n1971) );
  OAI21 U2087 ( .IN1(n714), .IN2(n1972), .IN3(n1971), .OUT(n1973) );
  AOI22 U2088 ( .IN1(n1974), .IN2(n1806), .IN3(RSTn), .IN4(n1973), .OUT(n1135)
         );
  MUX2X1 U2089 ( .IN1(n1983), .IN2(n1984), .S(n694), .OUT(n1554) );
  NOR2X1 U2090 ( .IN1(n695), .IN2(n694), .OUT(n1978) );
  INVX4 U2091 ( .IN(n1984), .OUT(n1981) );
  OAI21 U2092 ( .IN1(n695), .IN2(n1975), .IN3(n1981), .OUT(n1976) );
  OAI21 U2093 ( .IN1(n1978), .IN2(u_booth_count_reg_2_), .IN3(n1982), .OUT(
        n1980) );
  OAI21 U2094 ( .IN1(n1981), .IN2(n1980), .IN3(n1979), .OUT(n1555) );
  MUX2X1 U2095 ( .IN1(n1840), .IN2(u_booth_count_reg_3_), .S(n1982), .OUT(
        n1985) );
  AOI22 U2096 ( .IN1(n1985), .IN2(n1984), .IN3(u_booth_count_reg_3_), .IN4(
        n1983), .OUT(n1092) );
  NOR2X1 U2097 ( .IN1(n1986), .IN2(n2028), .OUT(n1987) );
  NOR2X1 U2098 ( .IN1(n715), .IN2(n1854), .OUT(Booth_dataout[1]) );
  NOR2X1 U2099 ( .IN1(n716), .IN2(n1786), .OUT(Booth_dataout[2]) );
  NOR2X1 U2100 ( .IN1(n718), .IN2(n1854), .OUT(Booth_dataout[4]) );
  NOR2X1 U2101 ( .IN1(n719), .IN2(n1854), .OUT(Booth_dataout[5]) );
  AOI22 U2102 ( .IN1(n2027), .IN2(MulCntrl_Op2[7]), .IN3(DIN2[7]), .IN4(n2026), 
        .OUT(n1992) );
  AOI22 U2103 ( .IN1(n2027), .IN2(n1862), .IN3(DIN2[8]), .IN4(n2026), .OUT(
        n1993) );
  AOI22 U2104 ( .IN1(n2027), .IN2(MulCntrl_Op2[9]), .IN3(DIN2[9]), .IN4(n2026), 
        .OUT(n1994) );
  AOI22 U2105 ( .IN1(n2027), .IN2(MulCntrl_Op2[10]), .IN3(DIN2[10]), .IN4(
        n2026), .OUT(n1995) );
  AOI22 U2106 ( .IN1(n2027), .IN2(MulCntrl_Op2[11]), .IN3(DIN2[11]), .IN4(
        n2026), .OUT(n1996) );
  AOI22 U2107 ( .IN1(n2027), .IN2(MulCntrl_Op2[12]), .IN3(DIN2[12]), .IN4(
        n2026), .OUT(n1997) );
  AOI22 U2108 ( .IN1(n2027), .IN2(n1863), .IN3(DIN2[13]), .IN4(n2026), .OUT(
        n1998) );
  AOI22 U2109 ( .IN1(n2027), .IN2(MulCntrl_Op2[14]), .IN3(DIN2[14]), .IN4(
        n2026), .OUT(n1999) );
  AOI22 U2110 ( .IN1(n2027), .IN2(MulCntrl_Op1[7]), .IN3(DIN1[7]), .IN4(n2026), 
        .OUT(n2000) );
  AOI22 U2111 ( .IN1(n2027), .IN2(n1865), .IN3(DIN1[8]), .IN4(n2026), .OUT(
        n2001) );
  AOI22 U2112 ( .IN1(n2027), .IN2(MulCntrl_Op1[9]), .IN3(DIN1[9]), .IN4(n2026), 
        .OUT(n2002) );
  AOI22 U2113 ( .IN1(n2027), .IN2(MulCntrl_Op1[10]), .IN3(DIN1[10]), .IN4(
        n2026), .OUT(n2003) );
  AOI22 U2114 ( .IN1(n2027), .IN2(MulCntrl_Op1[11]), .IN3(DIN1[11]), .IN4(
        n2026), .OUT(n2004) );
  AOI22 U2115 ( .IN1(n2027), .IN2(MulCntrl_Op1[12]), .IN3(DIN1[12]), .IN4(
        n2026), .OUT(n2005) );
  AOI22 U2116 ( .IN1(n2027), .IN2(MulCntrl_Op1[14]), .IN3(DIN1[14]), .IN4(
        n2026), .OUT(n2006) );
  AOI22 U2117 ( .IN1(Add_carryout), .IN2(n2008), .IN3(n2030), .IN4(
        u_adder_24b_N131), .OUT(n2007) );
  AOI22 U2118 ( .IN1(Add_dataout[7]), .IN2(n2008), .IN3(n2030), .IN4(
        u_adder_24b_N129), .OUT(n2009) );
  AOI22 U2119 ( .IN1(AdderCntrl_Op2[7]), .IN2(n2025), .IN3(DIN2[7]), .IN4(
        n1876), .OUT(n2013) );
  AOI22 U2120 ( .IN1(n2025), .IN2(n1870), .IN3(DIN2[8]), .IN4(n1876), .OUT(
        n2014) );
  AOI22 U2121 ( .IN1(n2025), .IN2(AdderCntrl_Op2[9]), .IN3(DIN2[9]), .IN4(
        n1876), .OUT(n2015) );
  AOI22 U2122 ( .IN1(n2025), .IN2(AdderCntrl_Op1[7]), .IN3(DIN1[7]), .IN4(
        n1876), .OUT(n2016) );
  AOI22 U2123 ( .IN1(n2025), .IN2(n1871), .IN3(DIN1[8]), .IN4(n1876), .OUT(
        n2017) );
  AOI22 U2124 ( .IN1(n2025), .IN2(n1869), .IN3(DIN1[9]), .IN4(n1876), .OUT(
        n2018) );
  AOI22 U2125 ( .IN1(n2022), .IN2(Add_dataout[6]), .IN3(n2021), .IN4(n1851), 
        .OUT(n2149) );
  AOI22 U2126 ( .IN1(n2022), .IN2(Add_dataout[7]), .IN3(n2021), .IN4(
        u_booth_A_reg_7_), .OUT(n2151) );
  AOI21 U2127 ( .IN1(u_booth_A_reg_7_), .IN2(n2024), .IN3(n709), .OUT(n2152)
         );
  NOR2X1 U2128 ( .IN1(MODE[1]), .IN2(MODE[0]), .OUT(n2045) );
  NOR2X1 U2129 ( .IN1(n2045), .IN2(MODE[2]), .OUT(n2043) );
  NAND3X1 U2130 ( .IN1(getdataStat_reg[0]), .IN2(n463), .IN3(ABUSY), .OUT(
        n2034) );
  NOR2X1 U2131 ( .IN1(n2034), .IN2(n1815), .OUT(AdderCntrl_valid) );
  NOR2X1 U2132 ( .IN1(ABUSY), .IN2(OPT), .OUT(n2035) );
  NAND3X1 U2133 ( .IN1(CS), .IN2(DIV), .IN3(n2035), .OUT(n2036) );
  NOR2X1 U2134 ( .IN1(getdataStat_reg[0]), .IN2(n2036), .OUT(n2221) );
  NOR2X1 U2135 ( .IN1(MBUSY), .IN2(getdataStat_reg[1]), .OUT(n2037) );
  NAND3X1 U2136 ( .IN1(DIV), .IN2(OPT), .IN3(n2037), .OUT(n2038) );
  NOR2X1 U2137 ( .IN1(n2086), .IN2(n2038), .OUT(n2204) );
  NOR2X1 U2138 ( .IN1(n2221), .IN2(n2204), .OUT(n2039) );
  INVX1 U2139 ( .IN(MODE[2]), .OUT(n2042) );
  AOI22 U2140 ( .IN1(MODE[2]), .IN2(n1817), .IN3(n463), .IN4(n2042), .OUT(
        n2040) );
  AOI22 U2141 ( .IN1(n2045), .IN2(n2040), .IN3(n2043), .IN4(
        AdderCntrl_Debug[0]), .OUT(n2041) );
  AOI22 U2142 ( .IN1(MODE[2]), .IN2(n1807), .IN3(n462), .IN4(n2042), .OUT(
        n2044) );
  AOI22 U2143 ( .IN1(n2045), .IN2(n2044), .IN3(n2043), .IN4(
        AdderCntrl_Debug[1]), .OUT(n2046) );
  NOR2X1 U2144 ( .IN1(n584), .IN2(n2078), .OUT(n2080) );
  NOR2X1 U2145 ( .IN1(n587), .IN2(n2086), .OUT(n2066) );
  AOI22 U2146 ( .IN1(n1872), .IN2(MultResult_reg[0]), .IN3(AdderResult_reg[0]), 
        .IN4(n1873), .OUT(n2047) );
  AOI22 U2147 ( .IN1(n1872), .IN2(MultResult_reg[10]), .IN3(
        AdderResult_reg[10]), .IN4(n1873), .OUT(n2048) );
  AOI22 U2148 ( .IN1(n1872), .IN2(MultResult_reg[11]), .IN3(
        AdderResult_reg[11]), .IN4(n1873), .OUT(n2049) );
  AOI22 U2149 ( .IN1(n1872), .IN2(MultResult_reg[12]), .IN3(
        AdderResult_reg[12]), .IN4(n1873), .OUT(n2050) );
  AOI22 U2150 ( .IN1(n1872), .IN2(MultResult_reg[13]), .IN3(
        AdderResult_reg[13]), .IN4(n1873), .OUT(n2051) );
  AOI22 U2151 ( .IN1(n1872), .IN2(MultResult_reg[14]), .IN3(
        AdderResult_reg[14]), .IN4(n1873), .OUT(n2052) );
  AOI22 U2152 ( .IN1(n1872), .IN2(MultResult_reg[15]), .IN3(
        AdderResult_reg[15]), .IN4(n1873), .OUT(n2053) );
  AOI22 U2153 ( .IN1(n1872), .IN2(MultResult_reg[1]), .IN3(AdderResult_reg[1]), 
        .IN4(n1873), .OUT(n2054) );
  AOI22 U2154 ( .IN1(n1872), .IN2(MultResult_reg[2]), .IN3(AdderResult_reg[2]), 
        .IN4(n1873), .OUT(n2055) );
  AOI22 U2155 ( .IN1(n1872), .IN2(MultResult_reg[3]), .IN3(AdderResult_reg[3]), 
        .IN4(n1873), .OUT(n2056) );
  AOI22 U2156 ( .IN1(n1872), .IN2(MultResult_reg[4]), .IN3(AdderResult_reg[4]), 
        .IN4(n1873), .OUT(n2057) );
  AOI22 U2157 ( .IN1(n1872), .IN2(MultResult_reg[5]), .IN3(AdderResult_reg[5]), 
        .IN4(n1873), .OUT(n2058) );
  AOI22 U2158 ( .IN1(n1872), .IN2(MultResult_reg[6]), .IN3(AdderResult_reg[6]), 
        .IN4(n1873), .OUT(n2059) );
  AOI22 U2159 ( .IN1(n1872), .IN2(MultResult_reg[7]), .IN3(AdderResult_reg[7]), 
        .IN4(n1873), .OUT(n2060) );
  AOI22 U2160 ( .IN1(n1872), .IN2(MultResult_reg[8]), .IN3(AdderResult_reg[8]), 
        .IN4(n1873), .OUT(n2061) );
  AOI22 U2161 ( .IN1(n1872), .IN2(MultResult_reg[9]), .IN3(AdderResult_reg[9]), 
        .IN4(n1873), .OUT(n2062) );
  NOR2X1 U2162 ( .IN1(n1872), .IN2(n1873), .OUT(n2063) );
  AOI22 U2163 ( .IN1(n1872), .IN2(MultExc_reg[0]), .IN3(AddExc_reg[0]), .IN4(
        n1873), .OUT(n2064) );
  AOI22 U2164 ( .IN1(n1872), .IN2(MultExc_reg[1]), .IN3(AddExc_reg[1]), .IN4(
        n1873), .OUT(n2065) );
  AOI22 U2165 ( .IN1(n1872), .IN2(MultExc_reg[2]), .IN3(AddExc_reg[2]), .IN4(
        n1873), .OUT(n2067) );
  NAND3X1 U2166 ( .IN1(getdataStat_reg[1]), .IN2(MBUSY), .IN3(n1817), .OUT(
        n2068) );
  NOR2X1 U2167 ( .IN1(multStateMC[1]), .IN2(n2068), .OUT(MulCntrl_valid) );
  NAND3X1 U2168 ( .IN1(n463), .IN2(n587), .IN3(n1815), .OUT(n2071) );
  OAI21 U2169 ( .IN1(getdataStat_reg[0]), .IN2(n2221), .IN3(n2071), .OUT(n2069) );
  NOR2X1 U2170 ( .IN1(n1877), .IN2(n2069), .OUT(N147) );
  NAND3X1 U2171 ( .IN1(multStateMC[1]), .IN2(n584), .IN3(n1817), .OUT(n2073)
         );
  OAI21 U2172 ( .IN1(getdataStat_reg[1]), .IN2(n2204), .IN3(n2073), .OUT(n2070) );
  NOR2X1 U2173 ( .IN1(n1877), .IN2(n2070), .OUT(N148) );
  NOR2X1 U2174 ( .IN1(n1815), .IN2(n463), .OUT(n2085) );
  INVX1 U2175 ( .IN(n2085), .OUT(n2075) );
  OAI21 U2176 ( .IN1(ABUSY), .IN2(n2221), .IN3(n2071), .OUT(n2072) );
  AOI21 U2177 ( .IN1(n2075), .IN2(n2072), .IN3(n1877), .OUT(N149) );
  OAI21 U2178 ( .IN1(MBUSY), .IN2(n2204), .IN3(n2073), .OUT(n2074) );
  AOI21 U2179 ( .IN1(n2156), .IN2(n2074), .IN3(n1877), .OUT(N150) );
  NOR2X1 U2180 ( .IN1(AdderCntrl_Dataout_valid), .IN2(n2075), .OUT(n2271) );
  NOR2X1 U2181 ( .IN1(n587), .IN2(n1877), .OUT(n2076) );
  OAI21 U2182 ( .IN1(n2270), .IN2(n2078), .IN3(n2077), .OUT(N189) );
  NAND2X1 U2183 ( .IN1(n1878), .IN2(n1848), .OUT(n2081) );
  NOR2X1 U2184 ( .IN1(n2156), .IN2(n2079), .OUT(n2248) );
  AOI21 U2185 ( .IN1(n2081), .IN2(n2155), .IN3(n1872), .OUT(N190) );
  NAND2X1 U2186 ( .IN1(n2082), .IN2(n2270), .OUT(N191) );
  AOI21 U2187 ( .IN1(n587), .IN2(n463), .IN3(n1877), .OUT(n2083) );
  NAND2X1 U2188 ( .IN1(n1815), .IN2(n2083), .OUT(n2084) );
  OAI21 U2189 ( .IN1(n2270), .IN2(n2086), .IN3(n2084), .OUT(n1692) );
  OAI21 U2190 ( .IN1(n2086), .IN2(AdderCntrl_Dataout_valid), .IN3(n2085), 
        .OUT(n2087) );
  NOR2X1 U2191 ( .IN1(AdderCntrl_valid), .IN2(n2088), .OUT(n2089) );
  OAI21 U2192 ( .IN1(n463), .IN2(n462), .IN3(n2089), .OUT(n2090) );
  NOR2X1 U2193 ( .IN1(u_ExcChecker_interconnect_stateMC_0_), .IN2(
        u_ExcChecker_interconnect_stateMC_1_), .OUT(n2103) );
  NAND2X1 U2194 ( .IN1(AdderCntrl_ExcCheck_valid), .IN2(n1825), .OUT(n2091) );
  AOI22 U2195 ( .IN1(u_ExcChecker_interconnect_stateMC_1_), .IN2(n1823), .IN3(
        n2103), .IN4(n2091), .OUT(n2093) );
  NAND2X1 U2196 ( .IN1(MulCntrl_ExcCheck_valid), .IN2(n1878), .OUT(n2092) );
  NAND3X1 U2197 ( .IN1(n1878), .IN2(u_ExcChecker_interconnect_stateMC_0_), 
        .IN3(u_ExcChecker_interconnect_stateMC_1_), .OUT(n2095) );
  OAI21 U2198 ( .IN1(n2093), .IN2(n2092), .IN3(n2095), .OUT(n1661) );
  NAND2X1 U2199 ( .IN1(MulCntrl_ExcCheck_valid), .IN2(
        u_ExcChecker_interconnect_priority_reg), .OUT(n2094) );
  AOI22 U2200 ( .IN1(u_ExcChecker_interconnect_stateMC_0_), .IN2(n1823), .IN3(
        n2103), .IN4(n2094), .OUT(n2097) );
  NAND2X1 U2201 ( .IN1(AdderCntrl_ExcCheck_valid), .IN2(n1878), .OUT(n2096) );
  OAI21 U2202 ( .IN1(n2097), .IN2(n2096), .IN3(n2095), .OUT(n1660) );
  INVX1 U2203 ( .IN(MulCntrl_ExcCheck_valid), .OUT(n2098) );
  AOI22 U2204 ( .IN1(u_ExcChecker_interconnect_priority_reg), .IN2(n2098), 
        .IN3(AdderCntrl_ExcCheck_valid), .IN4(n1825), .OUT(n2100) );
  OAI21 U2205 ( .IN1(u_ExcChecker_interconnect_priority_reg), .IN2(n2103), 
        .IN3(n1878), .OUT(n2099) );
  AOI21 U2206 ( .IN1(n2103), .IN2(n2100), .IN3(n2099), .OUT(n1659) );
  NAND3X1 U2207 ( .IN1(u_ExcChecker_interconnect_stateMC_1_), .IN2(
        MulCntrl_ExcCheck_valid), .IN3(n1820), .OUT(n2161) );
  NAND3X1 U2208 ( .IN1(u_ExcChecker_interconnect_stateMC_0_), .IN2(
        AdderCntrl_ExcCheck_valid), .IN3(n1827), .OUT(n2192) );
  NAND2X1 U2209 ( .IN1(ExcSelect), .IN2(n2192), .OUT(n2101) );
  AOI21 U2210 ( .IN1(n2161), .IN2(n2101), .IN3(n1877), .OUT(n1658) );
  AOI21 U2211 ( .IN1(ExcCheck_valid), .IN2(n1850), .IN3(u_exc_check_StateMC_0_), .OUT(n2102) );
  NOR2X1 U2212 ( .IN1(n2102), .IN2(n1877), .OUT(n1657) );
  NAND3X1 U2213 ( .IN1(n654), .IN2(ExcCheck_valid), .IN3(n1837), .OUT(n2106)
         );
  NOR2X1 U2214 ( .IN1(n1877), .IN2(n2106), .OUT(u_exc_check_N45) );
  NOR2X1 U2215 ( .IN1(n2103), .IN2(n1877), .OUT(n2195) );
  NOR2X1 U2216 ( .IN1(n1877), .IN2(n1823), .OUT(n2193) );
  AOI22 U2217 ( .IN1(n2195), .IN2(MulCntrl_Exc_Ack), .IN3(n2104), .IN4(n2193), 
        .OUT(n2105) );
  NOR2X1 U2218 ( .IN1(AdderCntrl_ExcCheck_Datain[3]), .IN2(
        AdderCntrl_ExcCheck_Datain[4]), .OUT(n2108) );
  NOR2X1 U2219 ( .IN1(AdderCntrl_ExcCheck_Datain[2]), .IN2(
        AdderCntrl_ExcCheck_Datain[0]), .OUT(n2107) );
  NOR2X1 U2220 ( .IN1(AdderCntrl_ExcCheck_Datain[1]), .IN2(n2109), .OUT(n2111)
         );
  NOR2X1 U2221 ( .IN1(AdderCntrl_ExcCheck_Datain[5]), .IN2(
        AdderCntrl_ExcCheck_Datain[6]), .OUT(n2110) );
  NAND3X1 U2222 ( .IN1(n2111), .IN2(n2110), .IN3(n1821), .OUT(n2122) );
  NOR2X1 U2223 ( .IN1(MulCntrl_ExcCheck_Datain[3]), .IN2(
        MulCntrl_ExcCheck_Datain[4]), .OUT(n2113) );
  NOR2X1 U2224 ( .IN1(MulCntrl_ExcCheck_Datain[2]), .IN2(
        MulCntrl_ExcCheck_Datain[0]), .OUT(n2112) );
  NOR2X1 U2225 ( .IN1(MulCntrl_ExcCheck_Datain[1]), .IN2(n2114), .OUT(n2116)
         );
  NOR2X1 U2226 ( .IN1(MulCntrl_ExcCheck_Datain[5]), .IN2(
        MulCntrl_ExcCheck_Datain[6]), .OUT(n2115) );
  NAND3X1 U2227 ( .IN1(n2116), .IN2(n2115), .IN3(ExcSelect), .OUT(n2127) );
  NOR2X1 U2228 ( .IN1(AdderCntrl_ExcCheck_Datain[14]), .IN2(
        AdderCntrl_ExcCheck_Datain[9]), .OUT(n2131) );
  INVX1 U2229 ( .IN(AdderCntrl_ExcCheck_Datain[13]), .OUT(n2117) );
  NOR2X1 U2230 ( .IN1(AdderCntrl_ExcCheck_Datain[12]), .IN2(n2117), .OUT(n2120) );
  NOR2X1 U2231 ( .IN1(AdderCntrl_ExcCheck_Datain[11]), .IN2(n1781), .OUT(n2119) );
  NOR2X1 U2232 ( .IN1(AdderCntrl_ExcCheck_Datain[8]), .IN2(n1782), .OUT(n2118)
         );
  NAND3X1 U2233 ( .IN1(n2120), .IN2(n2119), .IN3(n2118), .OUT(n2121) );
  NOR2X1 U2234 ( .IN1(n2122), .IN2(n2121), .OUT(n2130) );
  NOR2X1 U2235 ( .IN1(MulCntrl_ExcCheck_Datain[9]), .IN2(
        MulCntrl_ExcCheck_Datain[8]), .OUT(n2129) );
  NOR2X1 U2236 ( .IN1(MulCntrl_ExcCheck_Datain[12]), .IN2(
        MulCntrl_ExcCheck_Datain[11]), .OUT(n2125) );
  NOR2X1 U2237 ( .IN1(MulCntrl_ExcCheck_Datain[14]), .IN2(
        MulCntrl_ExcCheck_Datain[13]), .OUT(n2124) );
  NOR2X1 U2238 ( .IN1(MulCntrl_ExcCheck_Datain[7]), .IN2(
        MulCntrl_ExcCheck_Datain[10]), .OUT(n2123) );
  NAND3X1 U2239 ( .IN1(n2125), .IN2(n2124), .IN3(n2123), .OUT(n2126) );
  NOR2X1 U2240 ( .IN1(n2127), .IN2(n2126), .OUT(n2128) );
  AOI22 U2241 ( .IN1(n2131), .IN2(n2130), .IN3(n2129), .IN4(n2128), .OUT(n2197) );
  OAI21 U2242 ( .IN1(n2199), .IN2(n2132), .IN3(n2197), .OUT(n2133) );
  OAI21 U2243 ( .IN1(n2200), .IN2(n1824), .IN3(n2134), .OUT(n1655) );
  OAI21 U2244 ( .IN1(n2200), .IN2(n1847), .IN3(n2134), .OUT(n1654) );
  NOR2X1 U2245 ( .IN1(u_Adder_interconnect_stateMC_1_), .IN2(n1809), .OUT(
        n2145) );
  NAND2X1 U2246 ( .IN1(Add_valid), .IN2(n1826), .OUT(n2136) );
  AOI22 U2247 ( .IN1(u_Adder_interconnect_stateMC_1_), .IN2(n1838), .IN3(n2145), .IN4(n2136), .OUT(n2138) );
  NAND3X1 U2248 ( .IN1(n1878), .IN2(u_Adder_interconnect_stateMC_1_), .IN3(
        n1809), .OUT(n2140) );
  OAI21 U2249 ( .IN1(n2138), .IN2(n2137), .IN3(n2140), .OUT(n1622) );
  NAND2X1 U2250 ( .IN1(u_Adder_interconnect_priority_reg), .IN2(n1843), .OUT(
        n2139) );
  AOI22 U2251 ( .IN1(n2145), .IN2(n2139), .IN3(n1809), .IN4(n1838), .OUT(n2142) );
  NAND2X1 U2252 ( .IN1(n1878), .IN2(Add_valid), .OUT(n2141) );
  OAI21 U2253 ( .IN1(n2142), .IN2(n2141), .IN3(n2140), .OUT(n1621) );
  AOI22 U2254 ( .IN1(u_Adder_interconnect_priority_reg), .IN2(n692), .IN3(
        Add_valid), .IN4(n1826), .OUT(n2144) );
  OAI21 U2255 ( .IN1(u_Adder_interconnect_priority_reg), .IN2(n2145), .IN3(
        n1878), .OUT(n2143) );
  AOI21 U2256 ( .IN1(n2145), .IN2(n2144), .IN3(n2143), .OUT(n1620) );
  NOR2X1 U2257 ( .IN1(n1877), .IN2(n1838), .OUT(n2189) );
  NOR2X1 U2258 ( .IN1(n2145), .IN2(n1877), .OUT(n2188) );
  AOI22 U2259 ( .IN1(n2189), .IN2(n2146), .IN3(n2188), .IN4(n1846), .OUT(n2147) );
  NOR2X1 U2260 ( .IN1(n1877), .IN2(n1807), .OUT(n2153) );
  OAI21 U2261 ( .IN1(n1848), .IN2(multStateMC[0]), .IN3(n2153), .OUT(n2154) );
  NAND2X1 U2262 ( .IN1(n2155), .IN2(n2154), .OUT(n1513) );
  AOI21 U2263 ( .IN1(MulCntrl_Dataout_valid), .IN2(CS), .IN3(n2156), .OUT(
        n2157) );
  NOR2X1 U2264 ( .IN1(MulCntrl_valid), .IN2(n2157), .OUT(n2158) );
  OAI21 U2265 ( .IN1(n1807), .IN2(n1817), .IN3(n2158), .OUT(n2159) );
  NAND2X1 U2266 ( .IN1(n1823), .IN2(n1878), .OUT(n2160) );
  AOI21 U2267 ( .IN1(n2161), .IN2(n2192), .IN3(n2160), .OUT(
        u_ExcChecker_interconnect_N53) );
  NAND2X1 U2268 ( .IN1(n1814), .IN2(n1805), .OUT(n2176) );
  NOR2X1 U2269 ( .IN1(u_booth_M_reg_2_), .IN2(n2176), .OUT(n2172) );
  INVX1 U2270 ( .IN(n2172), .OUT(n2173) );
  NOR2X1 U2271 ( .IN1(n2173), .IN2(u_booth_M_reg_3_), .OUT(n2169) );
  INVX1 U2272 ( .IN(n2169), .OUT(n2170) );
  NOR2X1 U2273 ( .IN1(u_booth_M_reg_4_), .IN2(n2170), .OUT(n2166) );
  INVX1 U2274 ( .IN(n2166), .OUT(n2167) );
  NOR2X1 U2275 ( .IN1(n2167), .IN2(u_booth_M_reg_5_), .OUT(n2163) );
  INVX1 U2276 ( .IN(n2163), .OUT(n2164) );
  NOR2X1 U2277 ( .IN1(u_booth_M_reg_6_), .IN2(n2164), .OUT(n2162) );
  MUX2X1 U2278 ( .IN1(n2164), .IN2(n2163), .S(u_booth_M_reg_6_), .OUT(n2165)
         );
  MUX2X1 U2279 ( .IN1(n2167), .IN2(n2166), .S(u_booth_M_reg_5_), .OUT(n2168)
         );
  MUX2X1 U2280 ( .IN1(n2170), .IN2(n2169), .S(u_booth_M_reg_4_), .OUT(n2171)
         );
  MUX2X1 U2281 ( .IN1(n2173), .IN2(n2172), .S(u_booth_M_reg_3_), .OUT(n2174)
         );
  MUX2X1 U2282 ( .IN1(n2176), .IN2(n2175), .S(u_booth_M_reg_2_), .OUT(n2177)
         );
  NAND2X1 U2283 ( .IN1(u_exc_check_StateMC_0_), .IN2(n1878), .OUT(n2179) );
  INVX1 U2284 ( .IN(u_exc_check_N45), .OUT(n2178) );
  OAI21 U2285 ( .IN1(n654), .IN2(n2179), .IN3(n2178), .OUT(n622) );
  AOI22 U2286 ( .IN1(u_booth_M_reg_7_), .IN2(n2186), .IN3(n2028), .IN4(
        Booth_datain1[7]), .OUT(n2180) );
  AOI22 U2287 ( .IN1(u_booth_M_reg_6_), .IN2(n2186), .IN3(n2028), .IN4(
        Booth_datain1[6]), .OUT(n2181) );
  AOI22 U2288 ( .IN1(u_booth_M_reg_5_), .IN2(n2186), .IN3(n2028), .IN4(
        Booth_datain1[5]), .OUT(n2182) );
  AOI22 U2289 ( .IN1(u_booth_M_reg_4_), .IN2(n2186), .IN3(n2028), .IN4(
        Booth_datain1[4]), .OUT(n2183) );
  AOI22 U2290 ( .IN1(u_booth_M_reg_3_), .IN2(n2186), .IN3(n2028), .IN4(
        Booth_datain1[3]), .OUT(n2184) );
  AOI22 U2291 ( .IN1(u_booth_M_reg_2_), .IN2(n2186), .IN3(n2028), .IN4(
        Booth_datain1[2]), .OUT(n2185) );
  AOI22 U2292 ( .IN1(n2190), .IN2(n2189), .IN3(n2188), .IN4(Add_ack), .OUT(
        n2191) );
  AOI22 U2293 ( .IN1(n2195), .IN2(AdderCntrl_Exc_Ack), .IN3(n2194), .IN4(n2193), .OUT(n2196) );
  OAI21 U2294 ( .IN1(n2199), .IN2(n2198), .IN3(n2197), .OUT(n2202) );
  AOI22 U2295 ( .IN1(u_exc_check_N45), .IN2(n2202), .IN3(n2201), .IN4(
        ExcCheck_value[2]), .OUT(n2203) );
  AOI22 U2296 ( .IN1(DIN2[0]), .IN2(n2026), .IN3(n2027), .IN4(MulCntrl_Op2[0]), 
        .OUT(n2205) );
  AOI22 U2297 ( .IN1(n2027), .IN2(MulCntrl_Op2[1]), .IN3(n2026), .IN4(DIN2[1]), 
        .OUT(n2206) );
  AOI22 U2298 ( .IN1(n2027), .IN2(MulCntrl_Op2[2]), .IN3(n2026), .IN4(DIN2[2]), 
        .OUT(n2207) );
  AOI22 U2299 ( .IN1(n2027), .IN2(MulCntrl_Op2[3]), .IN3(n2026), .IN4(DIN2[3]), 
        .OUT(n2208) );
  AOI22 U2300 ( .IN1(n2027), .IN2(MulCntrl_Op2[4]), .IN3(n2026), .IN4(DIN2[4]), 
        .OUT(n2209) );
  AOI22 U2301 ( .IN1(n2027), .IN2(MulCntrl_Op2[5]), .IN3(n2026), .IN4(DIN2[5]), 
        .OUT(n2210) );
  AOI22 U2302 ( .IN1(n2027), .IN2(MulCntrl_Op2[6]), .IN3(n2026), .IN4(DIN2[6]), 
        .OUT(n2211) );
  AOI22 U2303 ( .IN1(n2027), .IN2(MulCntrl_Op2[15]), .IN3(n2026), .IN4(
        DIN2[15]), .OUT(n2212) );
  AOI22 U2304 ( .IN1(n2027), .IN2(MulCntrl_Op1[0]), .IN3(n2026), .IN4(DIN1[0]), 
        .OUT(n2213) );
  AOI22 U2305 ( .IN1(n2027), .IN2(MulCntrl_Op1[1]), .IN3(n2026), .IN4(DIN1[1]), 
        .OUT(n2214) );
  AOI22 U2306 ( .IN1(n2027), .IN2(MulCntrl_Op1[2]), .IN3(n2026), .IN4(DIN1[2]), 
        .OUT(n2215) );
  AOI22 U2307 ( .IN1(n2027), .IN2(MulCntrl_Op1[3]), .IN3(n2026), .IN4(DIN1[3]), 
        .OUT(n2216) );
  AOI22 U2308 ( .IN1(n2027), .IN2(MulCntrl_Op1[4]), .IN3(n2026), .IN4(DIN1[4]), 
        .OUT(n2217) );
  AOI22 U2309 ( .IN1(n2027), .IN2(MulCntrl_Op1[5]), .IN3(n2026), .IN4(DIN1[5]), 
        .OUT(n2218) );
  AOI22 U2310 ( .IN1(n2027), .IN2(MulCntrl_Op1[6]), .IN3(n2026), .IN4(DIN1[6]), 
        .OUT(n2219) );
  AOI22 U2311 ( .IN1(n2027), .IN2(MulCntrl_Op1[15]), .IN3(n2026), .IN4(
        DIN1[15]), .OUT(n2220) );
  AOI22 U2312 ( .IN1(DIN2[0]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op2[0]), .OUT(n2222) );
  AOI22 U2313 ( .IN1(DIN2[1]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op2[1]), .OUT(n2223) );
  AOI22 U2314 ( .IN1(DIN2[2]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op2[2]), .OUT(n2224) );
  AOI22 U2315 ( .IN1(DIN2[3]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op2[3]), .OUT(n2225) );
  AOI22 U2316 ( .IN1(DIN2[4]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op2[4]), .OUT(n2226) );
  AOI22 U2317 ( .IN1(DIN2[5]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op2[5]), .OUT(n2227) );
  AOI22 U2318 ( .IN1(DIN2[6]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op2[6]), .OUT(n2228) );
  AOI22 U2319 ( .IN1(DIN2[10]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op2[10]), .OUT(n2229) );
  AOI22 U2320 ( .IN1(DIN2[11]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op2[11]), .OUT(n2230) );
  AOI22 U2321 ( .IN1(DIN2[12]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op2[12]), .OUT(n2231) );
  AOI22 U2322 ( .IN1(DIN2[13]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op2[13]), .OUT(n2232) );
  AOI22 U2323 ( .IN1(DIN2[14]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op2[14]), .OUT(n2233) );
  AOI22 U2324 ( .IN1(DIN2[15]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op2[15]), .OUT(n2234) );
  AOI22 U2325 ( .IN1(DIN1[0]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op1[0]), .OUT(n2235) );
  AOI22 U2326 ( .IN1(DIN1[1]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op1[1]), .OUT(n2236) );
  AOI22 U2327 ( .IN1(DIN1[2]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op1[2]), .OUT(n2237) );
  AOI22 U2328 ( .IN1(DIN1[3]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op1[3]), .OUT(n2238) );
  AOI22 U2329 ( .IN1(DIN1[4]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op1[4]), .OUT(n2239) );
  AOI22 U2330 ( .IN1(DIN1[5]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op1[5]), .OUT(n2240) );
  AOI22 U2331 ( .IN1(DIN1[6]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op1[6]), .OUT(n2241) );
  AOI22 U2332 ( .IN1(DIN1[10]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op1[10]), .OUT(n2242) );
  AOI22 U2333 ( .IN1(DIN1[11]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op1[11]), .OUT(n2243) );
  AOI22 U2334 ( .IN1(DIN1[12]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op1[12]), .OUT(n2244) );
  AOI22 U2335 ( .IN1(DIN1[13]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op1[13]), .OUT(n2245) );
  AOI22 U2336 ( .IN1(DIN1[14]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op1[14]), .OUT(n2246) );
  AOI22 U2337 ( .IN1(DIN1[15]), .IN2(n1876), .IN3(n2025), .IN4(
        AdderCntrl_Op1[15]), .OUT(n2247) );
  NOR2X1 U2338 ( .IN1(n2248), .IN2(n1877), .OUT(n2267) );
  AOI22 U2339 ( .IN1(n2268), .IN2(MulCntrl_Dataout[15]), .IN3(n1874), .IN4(
        MultResult_reg[15]), .OUT(n2249) );
  AOI22 U2340 ( .IN1(n2268), .IN2(MulCntrl_Dataout[14]), .IN3(n1874), .IN4(
        MultResult_reg[14]), .OUT(n2250) );
  AOI22 U2341 ( .IN1(n2268), .IN2(MulCntrl_Dataout[13]), .IN3(n1874), .IN4(
        MultResult_reg[13]), .OUT(n2251) );
  AOI22 U2342 ( .IN1(n2268), .IN2(MulCntrl_Dataout[12]), .IN3(n1874), .IN4(
        MultResult_reg[12]), .OUT(n2252) );
  AOI22 U2343 ( .IN1(n2268), .IN2(MulCntrl_Dataout[11]), .IN3(n1874), .IN4(
        MultResult_reg[11]), .OUT(n2253) );
  AOI22 U2344 ( .IN1(n2268), .IN2(MulCntrl_Dataout[10]), .IN3(n1874), .IN4(
        MultResult_reg[10]), .OUT(n2254) );
  AOI22 U2345 ( .IN1(n2268), .IN2(MulCntrl_Dataout[9]), .IN3(n1874), .IN4(
        MultResult_reg[9]), .OUT(n2255) );
  AOI22 U2346 ( .IN1(n2268), .IN2(MulCntrl_Dataout[8]), .IN3(n1874), .IN4(
        MultResult_reg[8]), .OUT(n2256) );
  AOI22 U2347 ( .IN1(n2268), .IN2(MulCntrl_Dataout[7]), .IN3(n1874), .IN4(
        MultResult_reg[7]), .OUT(n2257) );
  AOI22 U2348 ( .IN1(n2268), .IN2(MulCntrl_Dataout[6]), .IN3(n1874), .IN4(
        MultResult_reg[6]), .OUT(n2258) );
  AOI22 U2349 ( .IN1(n2268), .IN2(MulCntrl_Dataout[5]), .IN3(n1874), .IN4(
        MultResult_reg[5]), .OUT(n2259) );
  AOI22 U2350 ( .IN1(n2268), .IN2(MulCntrl_Dataout[4]), .IN3(n1874), .IN4(
        MultResult_reg[4]), .OUT(n2260) );
  AOI22 U2351 ( .IN1(n2268), .IN2(MulCntrl_Dataout[3]), .IN3(n1874), .IN4(
        MultResult_reg[3]), .OUT(n2261) );
  AOI22 U2352 ( .IN1(n2268), .IN2(MulCntrl_Dataout[2]), .IN3(n1874), .IN4(
        MultResult_reg[2]), .OUT(n2262) );
  AOI22 U2353 ( .IN1(n2268), .IN2(MulCntrl_Dataout[1]), .IN3(n1874), .IN4(
        MultResult_reg[1]), .OUT(n2263) );
  AOI22 U2354 ( .IN1(n2268), .IN2(MulCntrl_Dataout[0]), .IN3(n1874), .IN4(
        MultResult_reg[0]), .OUT(n2264) );
  AOI22 U2355 ( .IN1(n2268), .IN2(MulCntrl_Exc[2]), .IN3(n1874), .IN4(
        MultExc_reg[2]), .OUT(n2265) );
  AOI22 U2356 ( .IN1(n2268), .IN2(MulCntrl_Exc[1]), .IN3(n1874), .IN4(
        MultExc_reg[1]), .OUT(n2266) );
  AOI22 U2357 ( .IN1(n2268), .IN2(MulCntrl_Exc[0]), .IN3(n1874), .IN4(
        MultExc_reg[0]), .OUT(n2269) );
  NOR2X1 U2358 ( .IN1(n2271), .IN2(n1877), .OUT(n2290) );
  AOI22 U2359 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[15]), .IN3(n1875), .IN4(
        AdderResult_reg[15]), .OUT(n2272) );
  AOI22 U2360 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[14]), .IN3(n1875), .IN4(
        AdderResult_reg[14]), .OUT(n2273) );
  AOI22 U2361 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[13]), .IN3(n1875), .IN4(
        AdderResult_reg[13]), .OUT(n2274) );
  AOI22 U2362 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[12]), .IN3(n1875), .IN4(
        AdderResult_reg[12]), .OUT(n2275) );
  AOI22 U2363 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[11]), .IN3(n1875), .IN4(
        AdderResult_reg[11]), .OUT(n2276) );
  AOI22 U2364 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[10]), .IN3(n1875), .IN4(
        AdderResult_reg[10]), .OUT(n2277) );
  AOI22 U2365 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[9]), .IN3(n1875), .IN4(
        AdderResult_reg[9]), .OUT(n2278) );
  AOI22 U2366 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[8]), .IN3(n1875), .IN4(
        AdderResult_reg[8]), .OUT(n2279) );
  AOI22 U2367 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[7]), .IN3(n1875), .IN4(
        AdderResult_reg[7]), .OUT(n2280) );
  AOI22 U2368 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[6]), .IN3(n1875), .IN4(
        AdderResult_reg[6]), .OUT(n2281) );
  AOI22 U2369 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[5]), .IN3(n1875), .IN4(
        AdderResult_reg[5]), .OUT(n2282) );
  AOI22 U2370 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[4]), .IN3(n1875), .IN4(
        AdderResult_reg[4]), .OUT(n2283) );
  AOI22 U2371 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[3]), .IN3(n1875), .IN4(
        AdderResult_reg[3]), .OUT(n2284) );
  AOI22 U2372 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[2]), .IN3(n1875), .IN4(
        AdderResult_reg[2]), .OUT(n2285) );
  AOI22 U2373 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[1]), .IN3(n1875), .IN4(
        AdderResult_reg[1]), .OUT(n2286) );
  AOI22 U2374 ( .IN1(n2291), .IN2(AdderCntrl_Dataout[0]), .IN3(n1875), .IN4(
        AdderResult_reg[0]), .OUT(n2287) );
  AOI22 U2375 ( .IN1(n2291), .IN2(AdderCntrl_Exc[2]), .IN3(n1875), .IN4(
        AddExc_reg[2]), .OUT(n2288) );
  AOI22 U2376 ( .IN1(n2291), .IN2(AdderCntrl_Exc[1]), .IN3(n1875), .IN4(
        AddExc_reg[1]), .OUT(n2289) );
  AOI22 U2377 ( .IN1(n2291), .IN2(AdderCntrl_Exc[0]), .IN3(n1875), .IN4(
        AddExc_reg[0]), .OUT(n2292) );
endmodule

