/home/arnabd/Semester1/DVLSI/Cadence-f15/Project/FPU/16edi_final/Lib6710_05.lef