
module Adder_cntrl ( CLK, RSTn, Datain1, Datain2, Data_valid, Dataout, Exc, 
        Mode, Debug, Adder_datain1, Adder_datain2, Adder_valid, Adder_dataout, 
        Adder_carryout, Adder_ack, ExcCheck_valid, Exc_value, Exc_Ack, 
        Dataout_valid_BAR, ExcCheck_Datain_15_, ExcCheck_Datain_14_, 
        ExcCheck_Datain_13__BAR, ExcCheck_Datain_12_, ExcCheck_Datain_11_, 
        ExcCheck_Datain_9_, ExcCheck_Datain_8_, ExcCheck_Datain_6_, 
        ExcCheck_Datain_5_, ExcCheck_Datain_4_, ExcCheck_Datain_3_, 
        ExcCheck_Datain_2_, ExcCheck_Datain_1_, ExcCheck_Datain_0_, 
        ExcCheck_Datain_10__BAR, ExcCheck_Datain_7__BAR );
  input [15:0] Datain1;
  input [15:0] Datain2;
  output [15:0] Dataout;
  output [2:0] Exc;
  input [2:0] Mode;
  output [4:0] Debug;
  output [8:0] Adder_datain1;
  output [8:0] Adder_datain2;
  input [8:0] Adder_dataout;
  input [2:0] Exc_value;
  input CLK, RSTn, Data_valid, Adder_carryout, Adder_ack, Exc_Ack;
  output Adder_valid, ExcCheck_valid, Dataout_valid_BAR, ExcCheck_Datain_15_,
         ExcCheck_Datain_14_, ExcCheck_Datain_13__BAR, ExcCheck_Datain_12_,
         ExcCheck_Datain_11_, ExcCheck_Datain_9_, ExcCheck_Datain_8_,
         ExcCheck_Datain_6_, ExcCheck_Datain_5_, ExcCheck_Datain_4_,
         ExcCheck_Datain_3_, ExcCheck_Datain_2_, ExcCheck_Datain_1_,
         ExcCheck_Datain_0_, ExcCheck_Datain_10__BAR, ExcCheck_Datain_7__BAR;
  wire   N148, N149, N150, N152, N156, N161, N162, N168, Debug_valid_reg,
         Op2_Mantissa_reg_7_, exc_reg_0_, carry_reg, N256, N257, N258, N259,
         N260, N261, N262, N263, N274, N366, N380, N434, N696, C493_DATA2_0,
         C493_DATA2_1, C493_DATA2_2, C493_DATA2_3, C493_DATA2_4, C493_DATA2_5,
         C493_DATA2_6, C493_DATA2_7, n73, n103, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n118, n119, n120, n121, n128, n191, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n217, n218, n274,
         n277, n665, n672, n958, n965, n1046, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         add_x_35_A_9_, add_x_35_A_8_, add_x_35_A_7_, add_x_35_A_6_,
         add_x_35_A_5_, add_x_35_A_4_, add_x_35_A_3_, add_x_35_A_2_,
         add_x_35_A_1_, add_x_35_A_0_, C1_Z_3, C1_Z_2, C1_Z_1, C1_Z_0, C2_Z_0,
         DP_OP_1074_157_5430_n34, DP_OP_1074_157_5430_n33,
         DP_OP_1074_157_5430_n32, DP_OP_1074_157_5430_n31,
         DP_OP_1074_157_5430_n30, DP_OP_1074_157_5430_n29,
         DP_OP_1074_157_5430_n28, DP_OP_1074_157_5430_n27,
         DP_OP_1074_157_5430_n26, DP_OP_1074_157_5430_n25,
         DP_OP_1074_157_5430_n24, DP_OP_1074_157_5430_n23,
         DP_OP_1074_157_5430_n22, DP_OP_1074_157_5430_n21,
         DP_OP_1074_157_5430_n20, DP_OP_1074_157_5430_n19,
         DP_OP_1074_157_5430_n14, DP_OP_1074_157_5430_n13,
         DP_OP_1074_157_5430_n12, DP_OP_1074_157_5430_n11,
         DP_OP_1074_157_5430_n10, DP_OP_1074_157_5430_n9,
         DP_OP_1074_157_5430_n8, DP_OP_1074_157_5430_n7,
         DP_OP_1074_157_5430_n6, DP_OP_1074_157_5430_n5,
         DP_OP_1074_157_5430_n4, DP_OP_1074_157_5430_n3,
         DP_OP_1074_157_5430_n2, DP_OP_1074_157_5430_n1, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n104, n115,
         n116, n117, n122, n123, n124, n125, n126, n127, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n216, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n275, n276,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n666, n667, n668, n669, n670, n671, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n822, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n959, n960, n961, n962, n963, n964,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225;
  wire   [2:0] StateMC;
  wire   [3:0] Debug_reg;
  wire   [7:0] Final_Exponent_reg;
  wire   [10:1] Final_Mantissa_reg;

  DFFRX1 Add_sign_reg_reg ( .D(n1165), .CLK(CLK), .CLRB(n73), .Q(n206), .QB(
        n277) );
  DFFRX1 StateMC_reg_1_ ( .D(n965), .CLK(CLK), .CLRB(n73), .Q(n199), .QB(
        StateMC[1]) );
  DFFRX1 Final_Mantissa_reg_reg_10_ ( .D(n1124), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[10]), .QB(n194) );
  DFFRX1 exc_reg_reg_0_ ( .D(n1154), .CLK(CLK), .CLRB(n73), .Q(exc_reg_0_), 
        .QB(n229) );
  DFFRX1 StateMC_reg_0_ ( .D(n1046), .CLK(CLK), .CLRB(n73), .Q(n223), .QB(
        StateMC[0]) );
  DFFRX1 StateMC_reg_2_ ( .D(n958), .CLK(CLK), .CLRB(n73), .Q(n198), .QB(
        StateMC[2]) );
  DFFRX1 Op2_Mantissa_reg_reg_6_ ( .D(n1136), .CLK(CLK), .CLRB(n73), .Q(n231), 
        .QB(add_x_35_A_9_) );
  DFFRX1 Op2_Mantissa_reg_reg_5_ ( .D(n1137), .CLK(CLK), .CLRB(n73), .Q(n228), 
        .QB(add_x_35_A_8_) );
  DFFRX1 Op2_Mantissa_reg_reg_4_ ( .D(n1138), .CLK(CLK), .CLRB(n73), .Q(n226), 
        .QB(add_x_35_A_7_) );
  DFFRX1 Op2_Mantissa_reg_reg_3_ ( .D(n1139), .CLK(CLK), .CLRB(n73), .Q(n225), 
        .QB(add_x_35_A_6_) );
  DFFRX1 Op2_Mantissa_reg_reg_2_ ( .D(n1140), .CLK(CLK), .CLRB(n73), .Q(n227), 
        .QB(add_x_35_A_5_) );
  DFFRX1 Op2_Mantissa_reg_reg_1_ ( .D(n1141), .CLK(CLK), .CLRB(n73), .Q(n232), 
        .QB(add_x_35_A_4_) );
  DFFRX1 Op2_Mantissa_reg_reg_0_ ( .D(n1142), .CLK(CLK), .CLRB(n73), .Q(n224), 
        .QB(add_x_35_A_3_) );
  DFFRX1 Op2_Mantissa_reg_reg_7_ ( .D(n1135), .CLK(CLK), .CLRB(n73), .Q(
        Op2_Mantissa_reg_7_), .QB(n239) );
  DFFRX1 exc_reg_reg_1_ ( .D(n1155), .CLK(CLK), .CLRB(n73), .Q(n236), .QB(n218) );
  DFFRX1 Adder_valid_reg ( .D(n1153), .CLK(CLK), .CLRB(n73), .Q(Adder_valid)
         );
  DFFRX1 Op1_Sign_reg_reg ( .D(n1143), .CLK(CLK), .CLRB(n73), .Q(n216), .QB(
        n191) );
  DFFRX1 Op1_Mantissa_reg_reg_6_ ( .D(n1145), .CLK(CLK), .CLRB(n73), .QB(n208)
         );
  DFFRX1 Adder_datain1_reg_6_ ( .D(N262), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[6]) );
  DFFRX1 Op1_Mantissa_reg_reg_5_ ( .D(n1146), .CLK(CLK), .CLRB(n73), .QB(n209)
         );
  DFFRX1 Adder_datain1_reg_5_ ( .D(N261), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[5]) );
  DFFRX1 Op1_Mantissa_reg_reg_4_ ( .D(n1147), .CLK(CLK), .CLRB(n73), .QB(n210)
         );
  DFFRX1 Adder_datain1_reg_4_ ( .D(N260), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[4]) );
  DFFRX1 Op1_Mantissa_reg_reg_3_ ( .D(n1148), .CLK(CLK), .CLRB(n73), .QB(n211)
         );
  DFFRX1 Adder_datain1_reg_3_ ( .D(N259), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[3]) );
  DFFRX1 Op1_Mantissa_reg_reg_2_ ( .D(n1149), .CLK(CLK), .CLRB(n73), .QB(n212)
         );
  DFFRX1 Adder_datain1_reg_2_ ( .D(N258), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[2]) );
  DFFRX1 Op1_Mantissa_reg_reg_1_ ( .D(n1150), .CLK(CLK), .CLRB(n73), .QB(n213)
         );
  DFFRX1 Adder_datain1_reg_1_ ( .D(N257), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[1]) );
  DFFRX1 Op1_Mantissa_reg_reg_0_ ( .D(n1151), .CLK(CLK), .CLRB(n73), .QB(n214)
         );
  DFFRX1 Adder_datain1_reg_0_ ( .D(N256), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[0]) );
  DFFRX1 Op2_Sign_reg_reg ( .D(n1152), .CLK(CLK), .CLRB(n73), .QB(n215) );
  DFFRX1 Adder_datain2_reg_8_ ( .D(n114), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[8]) );
  DFFRX1 Adder_datain2_reg_7_ ( .D(n113), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[7]) );
  DFFRX1 Adder_datain2_reg_6_ ( .D(n112), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[6]) );
  DFFRX1 Adder_datain2_reg_5_ ( .D(n111), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[5]) );
  DFFRX1 Adder_datain2_reg_4_ ( .D(n110), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[4]) );
  DFFRX1 Adder_datain2_reg_3_ ( .D(n109), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[3]) );
  DFFRX1 Adder_datain2_reg_2_ ( .D(n108), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[2]) );
  DFFRX1 Adder_datain2_reg_1_ ( .D(n107), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[1]) );
  DFFRX1 Adder_datain2_reg_0_ ( .D(n106), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[0]) );
  DFFRX1 R_reg_reg ( .D(n1132), .CLK(CLK), .CLRB(n73), .Q(n238), .QB(
        add_x_35_A_1_) );
  DFFRX1 S_reg_reg ( .D(n1133), .CLK(CLK), .CLRB(n73), .Q(n200), .QB(
        add_x_35_A_0_) );
  DFFRX1 G_reg_reg ( .D(n1134), .CLK(CLK), .CLRB(n73), .Q(n237), .QB(
        add_x_35_A_2_) );
  DFFRX1 Final_Mantissa_reg_reg_2_ ( .D(n665), .CLK(CLK), .CLRB(n73), .Q(n190), 
        .QB(Final_Mantissa_reg[2]) );
  DFFRX1 Final_Mantissa_reg_reg_1_ ( .D(n672), .CLK(CLK), .CLRB(n73), .Q(n192), 
        .QB(Final_Mantissa_reg[1]) );
  DFFRX1 Final_Mantissa_reg_reg_0_ ( .D(n128), .CLK(CLK), .CLRB(n73), .Q(N696), 
        .QB(n197) );
  DFFRX1 Final_Mantissa_reg_reg_8_ ( .D(n1126), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[8]), .QB(n195) );
  DFFRX1 Final_Mantissa_reg_reg_9_ ( .D(n1125), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[9]), .QB(n219) );
  DFFRX1 Final_Mantissa_reg_reg_7_ ( .D(n1127), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[7]), .QB(n204) );
  DFFRX1 Final_Mantissa_reg_reg_6_ ( .D(n1128), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[6]), .QB(n222) );
  DFFRX1 Final_Mantissa_reg_reg_5_ ( .D(n1129), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[5]), .QB(n193) );
  DFFRX1 Final_Mantissa_reg_reg_4_ ( .D(n1130), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[4]), .QB(n203) );
  DFFRX1 Final_Mantissa_reg_reg_3_ ( .D(n1131), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[3]), .QB(n201) );
  DFFRX1 carry_reg_reg ( .D(n1123), .CLK(CLK), .CLRB(n73), .Q(carry_reg), .QB(
        n221) );
  DFFRX1 Final_Exponent_reg_reg_0_ ( .D(n1156), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[0]), .QB(n220) );
  DFFRX1 Final_Exponent_reg_reg_1_ ( .D(n1157), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[1]), .QB(n196) );
  DFFRX1 Final_Exponent_reg_reg_2_ ( .D(n1158), .CLK(CLK), .CLRB(n73), .QB(
        n205) );
  DFFRX1 Final_Exponent_reg_reg_3_ ( .D(n1159), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[3]), .QB(n202) );
  DFFRX1 Final_Exponent_reg_reg_4_ ( .D(n1160), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[4]), .QB(n230) );
  DFFRX1 Final_Exponent_reg_reg_5_ ( .D(n1161), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[5]), .QB(n233) );
  DFFRX1 Final_Exponent_reg_reg_6_ ( .D(n1162), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[6]), .QB(n234) );
  DFFRX1 Final_Exponent_reg_reg_7_ ( .D(n1164), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[7]), .QB(n235) );
  DFFRX1 exc_reg_reg_2_ ( .D(n1163), .CLK(CLK), .CLRB(n73), .QB(n217) );
  DFFRX1 Op1_Mantissa_reg_reg_7_ ( .D(n1144), .CLK(CLK), .CLRB(n73), .QB(n207)
         );
  DFFRX1 Adder_datain1_reg_7_ ( .D(N263), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[7]) );
  DFFRX1 Debug_valid_reg_reg ( .D(n103), .CLK(CLK), .CLRB(n73), .Q(
        Debug_valid_reg), .QB(n240) );
  DFFRX1 Final_Sign_reg_reg ( .D(n1122), .CLK(CLK), .CLRB(n73), .Q(n241), .QB(
        n274) );
  DFFRX1 ExcCheck_valid_reg ( .D(N274), .CLK(CLK), .CLRB(n73), .Q(
        ExcCheck_valid) );
  DFFRX1 Debug_reg_reg_3_ ( .D(n121), .CLK(CLK), .CLRB(n73), .Q(Debug_reg[3])
         );
  DFFRX1 Debug_reg_reg_2_ ( .D(n120), .CLK(CLK), .CLRB(n73), .Q(Debug_reg[2])
         );
  DFFRX1 Debug_reg_reg_1_ ( .D(n119), .CLK(CLK), .CLRB(n73), .Q(Debug_reg[1])
         );
  DFFRX1 Debug_reg_reg_0_ ( .D(n118), .CLK(CLK), .CLRB(n73), .Q(Debug_reg[0])
         );
  NAND2X1 DP_OP_1074_157_5430_U1 ( .IN1(DP_OP_1074_157_5430_n2), .IN2(
        DP_OP_1074_157_5430_n1), .OUT(C493_DATA2_7) );
  NANDX2 DP_OP_1074_157_5430_U27 ( .IN1(C2_Z_0), .IN2(DP_OP_1074_157_5430_n29), 
        .OUT(DP_OP_1074_157_5430_n27) );
  NAND2X1 DP_OP_1074_157_5430_U32 ( .IN1(C1_Z_0), .IN2(DP_OP_1074_157_5430_n33), .OUT(DP_OP_1074_157_5430_n32) );
  NANDX2 DP_OP_1074_157_5430_U28 ( .IN1(C1_Z_1), .IN2(DP_OP_1074_157_5430_n29), 
        .OUT(DP_OP_1074_157_5430_n28) );
  NANDX2 DP_OP_1074_157_5430_U29 ( .IN1(C1_Z_1), .IN2(C2_Z_0), .OUT(
        DP_OP_1074_157_5430_n29) );
  NANDX2 DP_OP_1074_157_5430_U24 ( .IN1(C1_Z_2), .IN2(DP_OP_1074_157_5430_n25), 
        .OUT(DP_OP_1074_157_5430_n24) );
  NANDX2 DP_OP_1074_157_5430_U25 ( .IN1(C1_Z_2), .IN2(C2_Z_0), .OUT(
        DP_OP_1074_157_5430_n25) );
  NANDX2 DP_OP_1074_157_5430_U2 ( .IN1(DP_OP_1074_157_5430_n7), .IN2(
        DP_OP_1074_157_5430_n3), .OUT(DP_OP_1074_157_5430_n1) );
  NANDX2 DP_OP_1074_157_5430_U5 ( .IN1(DP_OP_1074_157_5430_n5), .IN2(
        DP_OP_1074_157_5430_n4), .OUT(DP_OP_1074_157_5430_n7) );
  NANDX2 DP_OP_1074_157_5430_U30 ( .IN1(DP_OP_1074_157_5430_n32), .IN2(
        DP_OP_1074_157_5430_n31), .OUT(DP_OP_1074_157_5430_n34) );
  NANDX2 DP_OP_1074_157_5430_U26 ( .IN1(DP_OP_1074_157_5430_n28), .IN2(
        DP_OP_1074_157_5430_n27), .OUT(DP_OP_1074_157_5430_n30) );
  NANDX2 DP_OP_1074_157_5430_U22 ( .IN1(DP_OP_1074_157_5430_n24), .IN2(
        DP_OP_1074_157_5430_n23), .OUT(DP_OP_1074_157_5430_n26) );
  NANDX2 DP_OP_1074_157_5430_U18 ( .IN1(DP_OP_1074_157_5430_n20), .IN2(
        DP_OP_1074_157_5430_n19), .OUT(DP_OP_1074_157_5430_n22) );
  NANDX2 DP_OP_1074_157_5430_U20 ( .IN1(C1_Z_3), .IN2(DP_OP_1074_157_5430_n21), 
        .OUT(DP_OP_1074_157_5430_n20) );
  NANDX2 DP_OP_1074_157_5430_U21 ( .IN1(C1_Z_3), .IN2(C2_Z_0), .OUT(
        DP_OP_1074_157_5430_n21) );
  NAND2X1 DP_OP_1074_157_5430_U3 ( .IN1(DP_OP_1074_157_5430_n8), .IN2(
        DP_OP_1074_157_5430_n3), .OUT(DP_OP_1074_157_5430_n2) );
  NAND2X1 DP_OP_1074_157_5430_U4 ( .IN1(DP_OP_1074_157_5430_n8), .IN2(
        DP_OP_1074_157_5430_n7), .OUT(DP_OP_1074_157_5430_n3) );
  NAND2X1 DP_OP_1074_157_5430_U6 ( .IN1(Final_Exponent_reg[7]), .IN2(
        DP_OP_1074_157_5430_n6), .OUT(DP_OP_1074_157_5430_n4) );
  NAND2X1 DP_OP_1074_157_5430_U7 ( .IN1(C2_Z_0), .IN2(DP_OP_1074_157_5430_n6), 
        .OUT(DP_OP_1074_157_5430_n5) );
  NAND2X1 DP_OP_1074_157_5430_U8 ( .IN1(C2_Z_0), .IN2(Final_Exponent_reg[7]), 
        .OUT(DP_OP_1074_157_5430_n6) );
  FULLADD DP_OP_1074_157_5430_U15 ( .A(C2_Z_0), .B(n181), .CIN(
        DP_OP_1074_157_5430_n34), .COUT(DP_OP_1074_157_5430_n14), .SUM(
        C493_DATA2_0) );
  FULLADD DP_OP_1074_157_5430_U14 ( .A(DP_OP_1074_157_5430_n30), .B(
        Final_Exponent_reg[1]), .CIN(n176), .COUT(DP_OP_1074_157_5430_n13), 
        .SUM(C493_DATA2_1) );
  FULLADD DP_OP_1074_157_5430_U13 ( .A(DP_OP_1074_157_5430_n26), .B(n184), 
        .CIN(n187), .COUT(DP_OP_1074_157_5430_n12), .SUM(C493_DATA2_2) );
  FULLADD DP_OP_1074_157_5430_U12 ( .A(DP_OP_1074_157_5430_n22), .B(n183), 
        .CIN(n188), .COUT(DP_OP_1074_157_5430_n11), .SUM(C493_DATA2_3) );
  FULLADD DP_OP_1074_157_5430_U11 ( .A(C2_Z_0), .B(Final_Exponent_reg[4]), 
        .CIN(DP_OP_1074_157_5430_n11), .COUT(DP_OP_1074_157_5430_n10), .SUM(
        C493_DATA2_4) );
  FULLADD DP_OP_1074_157_5430_U10 ( .A(C2_Z_0), .B(n182), .CIN(n189), .COUT(
        DP_OP_1074_157_5430_n9), .SUM(C493_DATA2_5) );
  FULLADD DP_OP_1074_157_5430_U9 ( .A(C2_Z_0), .B(n180), .CIN(n178), .COUT(
        DP_OP_1074_157_5430_n8), .SUM(C493_DATA2_6) );
  NAND2X1 DP_OP_1074_157_5430_U33 ( .IN1(C1_Z_0), .IN2(C2_Z_0), .OUT(
        DP_OP_1074_157_5430_n33) );
  NAND2X1 DP_OP_1074_157_5430_U23 ( .IN1(C2_Z_0), .IN2(DP_OP_1074_157_5430_n25), .OUT(DP_OP_1074_157_5430_n23) );
  NAND2X1 DP_OP_1074_157_5430_U19 ( .IN1(C2_Z_0), .IN2(DP_OP_1074_157_5430_n21), .OUT(DP_OP_1074_157_5430_n19) );
  NAND3X1 U3 ( .IN1(n578), .IN2(n657), .IN3(n606), .OUT(n1) );
  INVX1 U4 ( .IN(n1), .OUT(n2) );
  NAND3X1 U5 ( .IN1(n644), .IN2(n587), .IN3(n2), .OUT(n681) );
  INVX1 U6 ( .IN(n1081), .OUT(n3) );
  OAI21 U7 ( .IN1(n363), .IN2(n3), .IN3(n1106), .OUT(n455) );
  INVX1 U8 ( .IN(n1193), .OUT(n4) );
  OAI21 U9 ( .IN1(n755), .IN2(n1086), .IN3(n696), .OUT(n5) );
  AOI22 U10 ( .IN1(Debug_reg[3]), .IN2(n1117), .IN3(n4), .IN4(n5), .OUT(n6) );
  INVX1 U11 ( .IN(n6), .OUT(n121) );
  NAND3X1 U12 ( .IN1(n261), .IN2(n195), .IN3(n714), .OUT(n657) );
  NAND2X1 U13 ( .IN1(n1190), .IN2(Debug_valid_reg), .OUT(n7) );
  NOR2X1 U14 ( .IN1(n724), .IN2(n723), .OUT(n8) );
  NAND3X1 U15 ( .IN1(n728), .IN2(n727), .IN3(n8), .OUT(n9) );
  NAND2X1 U16 ( .IN1(n725), .IN2(n726), .OUT(n10) );
  OAI21 U17 ( .IN1(n9), .IN2(n10), .IN3(n733), .OUT(n11) );
  OAI21 U18 ( .IN1(n732), .IN2(n731), .IN3(n1115), .OUT(n12) );
  NAND2X1 U19 ( .IN1(n12), .IN2(Mode[0]), .OUT(n13) );
  AOI21 U20 ( .IN1(n730), .IN2(n729), .IN3(n13), .OUT(n14) );
  NAND2X1 U21 ( .IN1(n11), .IN2(n14), .OUT(n15) );
  OAI21 U22 ( .IN1(n675), .IN2(n15), .IN3(n1192), .OUT(n16) );
  AOI22 U23 ( .IN1(n1193), .IN2(n7), .IN3(n240), .IN4(n16), .OUT(n103) );
  INVX1 U24 ( .IN(n1084), .OUT(n17) );
  AOI22 U25 ( .IN1(n517), .IN2(n262), .IN3(Final_Mantissa_reg[1]), .IN4(n750), 
        .OUT(n18) );
  INVX1 U26 ( .IN(n485), .OUT(n19) );
  AOI21 U27 ( .IN1(n360), .IN2(n193), .IN3(n19), .OUT(n20) );
  AOI22 U28 ( .IN1(n20), .IN2(n511), .IN3(Adder_dataout[2]), .IN4(n1088), 
        .OUT(n21) );
  OAI21 U29 ( .IN1(n222), .IN2(n512), .IN3(n21), .OUT(n22) );
  AOI21 U30 ( .IN1(n513), .IN2(n688), .IN3(n22), .OUT(n23) );
  OAI21 U31 ( .IN1(n382), .IN2(n18), .IN3(n23), .OUT(n24) );
  AOI21 U32 ( .IN1(n754), .IN2(n520), .IN3(n24), .OUT(n25) );
  OAI21 U33 ( .IN1(n482), .IN2(n17), .IN3(n25), .OUT(n26) );
  AOI21 U34 ( .IN1(n522), .IN2(n492), .IN3(n26), .OUT(n27) );
  NAND2X1 U35 ( .IN1(Final_Mantissa_reg[5]), .IN2(n490), .OUT(n28) );
  OAI21 U36 ( .IN1(n265), .IN2(n27), .IN3(n28), .OUT(n1129) );
  INVX1 U37 ( .IN(n531), .OUT(n29) );
  NOR2X1 U38 ( .IN1(n532), .IN2(n29), .OUT(n835) );
  AOI22 U39 ( .IN1(n258), .IN2(n487), .IN3(n260), .IN4(n750), .OUT(n30) );
  AOI22 U40 ( .IN1(Final_Mantissa_reg[5]), .IN2(n517), .IN3(n518), .IN4(n259), 
        .OUT(n31) );
  AOI21 U41 ( .IN1(n30), .IN2(n31), .IN3(n488), .OUT(n32) );
  AOI21 U42 ( .IN1(n222), .IN2(n485), .IN3(n484), .OUT(n33) );
  AOI22 U43 ( .IN1(n1088), .IN2(Adder_dataout[3]), .IN3(n33), .IN4(n511), 
        .OUT(n34) );
  OAI21 U44 ( .IN1(n204), .IN2(n512), .IN3(n34), .OUT(n35) );
  NOR2X1 U45 ( .IN1(n32), .IN2(n35), .OUT(n36) );
  AOI22 U46 ( .IN1(n524), .IN2(n513), .IN3(n521), .IN4(n486), .OUT(n37) );
  NAND2X1 U47 ( .IN1(n36), .IN2(n37), .OUT(n38) );
  AOI21 U48 ( .IN1(n522), .IN2(n489), .IN3(n38), .OUT(n39) );
  AOI22 U49 ( .IN1(n689), .IN2(n692), .IN3(n688), .IN4(n687), .OUT(n40) );
  AOI22 U50 ( .IN1(n524), .IN2(n751), .IN3(n691), .IN4(n686), .OUT(n41) );
  NAND2X1 U51 ( .IN1(n40), .IN2(n41), .OUT(n42) );
  AOI22 U52 ( .IN1(n260), .IN2(n490), .IN3(n527), .IN4(n42), .OUT(n43) );
  OAI21 U53 ( .IN1(n265), .IN2(n39), .IN3(n43), .OUT(n1128) );
  AOI22 U54 ( .IN1(n654), .IN2(n653), .IN3(n651), .IN4(n652), .OUT(n44) );
  INVX1 U55 ( .IN(n657), .OUT(n45) );
  AOI22 U56 ( .IN1(n660), .IN2(n45), .IN3(n659), .IN4(n658), .OUT(n46) );
  NOR2X1 U57 ( .IN1(n656), .IN2(n655), .OUT(n47) );
  NAND2X1 U58 ( .IN1(n44), .IN2(n46), .OUT(n48) );
  NOR2X1 U59 ( .IN1(n47), .IN2(n48), .OUT(n743) );
  NAND2X1 U60 ( .IN1(n264), .IN2(N168), .OUT(n49) );
  AOI21 U61 ( .IN1(n1067), .IN2(n49), .IN3(n1071), .OUT(n50) );
  INVX1 U62 ( .IN(n49), .OUT(n51) );
  AOI22 U63 ( .IN1(n51), .IN2(n929), .IN3(n992), .IN4(n49), .OUT(n52) );
  INVX1 U64 ( .IN(N156), .OUT(n53) );
  AOI22 U65 ( .IN1(N156), .IN2(n1203), .IN3(n1202), .IN4(n53), .OUT(n54) );
  AOI22 U66 ( .IN1(N156), .IN2(n1201), .IN3(n1200), .IN4(n53), .OUT(n55) );
  INVX1 U67 ( .IN(n52), .OUT(n56) );
  AOI22 U68 ( .IN1(n52), .IN2(n54), .IN3(n55), .IN4(n56), .OUT(n57) );
  AOI22 U69 ( .IN1(N156), .IN2(n1207), .IN3(n1206), .IN4(n53), .OUT(n58) );
  AOI22 U70 ( .IN1(N156), .IN2(n1205), .IN3(n1204), .IN4(n53), .OUT(n59) );
  AOI22 U71 ( .IN1(n52), .IN2(n58), .IN3(n59), .IN4(n56), .OUT(n60) );
  NAND2X1 U72 ( .IN1(n929), .IN2(n49), .OUT(n61) );
  MUX2X1 U73 ( .IN1(n772), .IN2(n913), .S(n61), .OUT(n62) );
  MUX2X1 U74 ( .IN1(n57), .IN2(n60), .S(n62), .OUT(n63) );
  NAND2X1 U75 ( .IN1(n1119), .IN2(n1068), .OUT(n64) );
  AOI22 U76 ( .IN1(n50), .IN2(n63), .IN3(n200), .IN4(n64), .OUT(n65) );
  INVX1 U77 ( .IN(N168), .OUT(n66) );
  AOI22 U78 ( .IN1(N168), .IN2(n1219), .IN3(n1218), .IN4(n66), .OUT(n67) );
  AOI22 U79 ( .IN1(N168), .IN2(n1221), .IN3(n1220), .IN4(n66), .OUT(n68) );
  NOR2X1 U80 ( .IN1(n179), .IN2(n984), .OUT(n69) );
  INVX1 U81 ( .IN(n1066), .OUT(n70) );
  AOI22 U82 ( .IN1(n69), .IN2(N156), .IN3(n984), .IN4(n70), .OUT(n71) );
  MUX2X1 U83 ( .IN1(n67), .IN2(n68), .S(n71), .OUT(n72) );
  AOI22 U84 ( .IN1(N168), .IN2(n1223), .IN3(n1222), .IN4(n66), .OUT(n74) );
  AOI22 U85 ( .IN1(N168), .IN2(n1225), .IN3(n1224), .IN4(n66), .OUT(n75) );
  MUX2X1 U86 ( .IN1(n74), .IN2(n75), .S(n71), .OUT(n76) );
  AOI21 U87 ( .IN1(N156), .IN2(N366), .IN3(n984), .OUT(n77) );
  MUX2X1 U88 ( .IN1(n893), .IN2(n784), .S(n77), .OUT(n78) );
  MUX2X1 U89 ( .IN1(n72), .IN2(n76), .S(n78), .OUT(n79) );
  NOR2X1 U90 ( .IN1(n1073), .IN2(n79), .OUT(n80) );
  OAI21 U91 ( .IN1(n1066), .IN2(n1065), .IN3(n80), .OUT(n81) );
  NAND2X1 U92 ( .IN1(n65), .IN2(n81), .OUT(n1133) );
  AOI22 U93 ( .IN1(n630), .IN2(n658), .IN3(n723), .IN4(n631), .OUT(n82) );
  INVX1 U94 ( .IN(n632), .OUT(n83) );
  NOR2X1 U95 ( .IN1(n708), .IN2(n633), .OUT(n84) );
  AOI21 U96 ( .IN1(n83), .IN2(n660), .IN3(n84), .OUT(n85) );
  NAND2X1 U97 ( .IN1(n82), .IN2(n85), .OUT(n86) );
  AOI21 U98 ( .IN1(n654), .IN2(n634), .IN3(n86), .OUT(n87) );
  OAI21 U99 ( .IN1(n635), .IN2(n725), .IN3(n87), .OUT(n88) );
  INVX1 U100 ( .IN(n636), .OUT(n89) );
  AOI22 U101 ( .IN1(n639), .IN2(n710), .IN3(n640), .IN4(n89), .OUT(n90) );
  OAI21 U102 ( .IN1(n628), .IN2(n643), .IN3(n90), .OUT(n91) );
  NOR2X1 U103 ( .IN1(n88), .IN2(n91), .OUT(n677) );
  NAND3X1 U104 ( .IN1(n180), .IN2(n182), .IN3(Final_Exponent_reg[7]), .OUT(n92) );
  INVX1 U105 ( .IN(n92), .OUT(n93) );
  INVX1 U106 ( .IN(n184), .OUT(n94) );
  NAND3X1 U107 ( .IN1(n183), .IN2(n181), .IN3(Final_Exponent_reg[1]), .OUT(n95) );
  NOR2X1 U108 ( .IN1(n94), .IN2(n95), .OUT(n96) );
  NAND3X1 U109 ( .IN1(Final_Exponent_reg[4]), .IN2(n93), .IN3(n96), .OUT(n532)
         );
  AOI22 U110 ( .IN1(Final_Mantissa_reg[8]), .IN2(n517), .IN3(n518), .IN4(n261), 
        .OUT(n97) );
  OAI21 U111 ( .IN1(n222), .IN2(n519), .IN3(n97), .OUT(n98) );
  AOI22 U112 ( .IN1(n520), .IN2(n521), .IN3(n754), .IN4(n98), .OUT(n99) );
  NOR2X1 U113 ( .IN1(Final_Mantissa_reg[9]), .IN2(n510), .OUT(n100) );
  AOI22 U114 ( .IN1(n511), .IN2(n100), .IN3(Adder_dataout[6]), .IN4(n1088), 
        .OUT(n101) );
  OAI21 U115 ( .IN1(n194), .IN2(n512), .IN3(n101), .OUT(n102) );
  AOI21 U116 ( .IN1(n525), .IN2(n513), .IN3(n102), .OUT(n104) );
  OAI21 U117 ( .IN1(n515), .IN2(n514), .IN3(n104), .OUT(n115) );
  AOI21 U118 ( .IN1(Final_Mantissa_reg[9]), .IN2(n516), .IN3(n115), .OUT(n116)
         );
  NAND2X1 U119 ( .IN1(n1084), .IN2(n522), .OUT(n117) );
  NAND3X1 U120 ( .IN1(n99), .IN2(n116), .IN3(n117), .OUT(n122) );
  NOR2X1 U121 ( .IN1(n509), .IN2(n508), .OUT(n123) );
  NOR2X1 U122 ( .IN1(n122), .IN2(n123), .OUT(n124) );
  AOI22 U123 ( .IN1(n525), .IN2(n751), .IN3(n526), .IN4(n691), .OUT(n125) );
  AOI22 U124 ( .IN1(n687), .IN2(n523), .IN3(n524), .IN4(n689), .OUT(n126) );
  NAND2X1 U125 ( .IN1(n125), .IN2(n126), .OUT(n127) );
  AOI22 U126 ( .IN1(Final_Mantissa_reg[9]), .IN2(n528), .IN3(n527), .IN4(n127), 
        .OUT(n129) );
  OAI21 U127 ( .IN1(n265), .IN2(n124), .IN3(n129), .OUT(n1125) );
  NOR2X1 U128 ( .IN1(n1072), .IN2(n1071), .OUT(n130) );
  INVX1 U129 ( .IN(N366), .OUT(n131) );
  AOI22 U130 ( .IN1(N366), .IN2(Datain2[3]), .IN3(Datain2[2]), .IN4(n131), 
        .OUT(n132) );
  AOI22 U131 ( .IN1(N366), .IN2(Datain2[1]), .IN3(Datain2[0]), .IN4(n131), 
        .OUT(n133) );
  INVX1 U132 ( .IN(n251), .OUT(n134) );
  AOI22 U133 ( .IN1(n251), .IN2(n132), .IN3(n133), .IN4(n134), .OUT(n135) );
  AOI22 U134 ( .IN1(N366), .IN2(Datain2[7]), .IN3(Datain2[6]), .IN4(n131), 
        .OUT(n136) );
  AOI22 U135 ( .IN1(N366), .IN2(Datain2[5]), .IN3(Datain2[4]), .IN4(n131), 
        .OUT(n137) );
  AOI22 U136 ( .IN1(n251), .IN2(n136), .IN3(n137), .IN4(n134), .OUT(n138) );
  AOI22 U137 ( .IN1(n929), .IN2(N168), .IN3(n251), .IN4(n992), .OUT(n139) );
  MUX2X1 U138 ( .IN1(n135), .IN2(n138), .S(n139), .OUT(n140) );
  AOI22 U139 ( .IN1(N366), .IN2(Datain2[11]), .IN3(Datain2[10]), .IN4(n131), 
        .OUT(n141) );
  INVX1 U140 ( .IN(n264), .OUT(n142) );
  AOI22 U141 ( .IN1(n264), .IN2(Datain2[9]), .IN3(Datain2[8]), .IN4(n142), 
        .OUT(n143) );
  AOI22 U142 ( .IN1(n251), .IN2(n141), .IN3(n143), .IN4(n134), .OUT(n144) );
  AOI22 U143 ( .IN1(n264), .IN2(Datain2[15]), .IN3(Datain2[14]), .IN4(n142), 
        .OUT(n145) );
  AOI22 U144 ( .IN1(N366), .IN2(Datain2[13]), .IN3(Datain2[12]), .IN4(n131), 
        .OUT(n146) );
  AOI22 U145 ( .IN1(n251), .IN2(n145), .IN3(n146), .IN4(n134), .OUT(n147) );
  MUX2X1 U146 ( .IN1(n144), .IN2(n147), .S(n139), .OUT(n148) );
  NOR2X1 U147 ( .IN1(N168), .IN2(n992), .OUT(n149) );
  MUX2X1 U148 ( .IN1(n913), .IN2(n772), .S(n149), .OUT(n150) );
  MUX2X1 U149 ( .IN1(n140), .IN2(n148), .S(n150), .OUT(n151) );
  AOI22 U150 ( .IN1(n997), .IN2(N156), .IN3(n252), .IN4(n984), .OUT(n152) );
  INVX1 U151 ( .IN(n252), .OUT(n153) );
  AOI22 U152 ( .IN1(n252), .IN2(n1217), .IN3(n1216), .IN4(n153), .OUT(n154) );
  AOI22 U153 ( .IN1(n252), .IN2(n1215), .IN3(n1214), .IN4(n153), .OUT(n155) );
  INVX1 U154 ( .IN(n152), .OUT(n156) );
  AOI22 U155 ( .IN1(n152), .IN2(n154), .IN3(n155), .IN4(n156), .OUT(n157) );
  AOI22 U156 ( .IN1(N366), .IN2(Datain1[11]), .IN3(Datain1[10]), .IN4(n131), 
        .OUT(n158) );
  AOI22 U157 ( .IN1(N366), .IN2(Datain1[9]), .IN3(Datain1[8]), .IN4(n131), 
        .OUT(n159) );
  AOI22 U158 ( .IN1(n252), .IN2(n158), .IN3(n159), .IN4(n153), .OUT(n160) );
  AOI22 U159 ( .IN1(N366), .IN2(Datain1[15]), .IN3(Datain1[14]), .IN4(n131), 
        .OUT(n161) );
  AOI22 U160 ( .IN1(N366), .IN2(Datain1[13]), .IN3(Datain1[12]), .IN4(n131), 
        .OUT(n162) );
  AOI22 U161 ( .IN1(n252), .IN2(n161), .IN3(n162), .IN4(n153), .OUT(n163) );
  MUX2X1 U162 ( .IN1(n160), .IN2(n163), .S(n152), .OUT(n164) );
  NOR2X1 U163 ( .IN1(N156), .IN2(n984), .OUT(n165) );
  AOI22 U164 ( .IN1(n893), .IN2(n984), .IN3(n784), .IN4(n165), .OUT(n166) );
  OAI21 U165 ( .IN1(n252), .IN2(n784), .IN3(n166), .OUT(n167) );
  MUX2X1 U166 ( .IN1(n157), .IN2(n164), .S(n167), .OUT(n168) );
  AOI21 U167 ( .IN1(n1075), .IN2(n1074), .IN3(n1073), .OUT(n169) );
  AOI22 U168 ( .IN1(n130), .IN2(n151), .IN3(n168), .IN4(n169), .OUT(n170) );
  MUX2X1 U169 ( .IN1(add_x_35_A_1_), .IN2(n238), .S(add_x_35_A_0_), .OUT(n171)
         );
  AOI22 U170 ( .IN1(n1069), .IN2(n238), .IN3(n1070), .IN4(n171), .OUT(n172) );
  NAND2X1 U171 ( .IN1(n170), .IN2(n172), .OUT(n1132) );
  INVX4 U172 ( .IN(n723), .OUT(n173) );
  NANDX2 U173 ( .IN1(Final_Mantissa_reg[10]), .IN2(n299), .OUT(n300) );
  NANDX2 U174 ( .IN1(n192), .IN2(n197), .OUT(n174) );
  INVX4 U175 ( .IN(n174), .OUT(n362) );
  INVX4 U176 ( .IN(n632), .OUT(n595) );
  NANDX2 U177 ( .IN1(n194), .IN2(n298), .OUT(n301) );
  INVX1 U178 ( .IN(DP_OP_1074_157_5430_n14), .OUT(n175) );
  INVX4 U179 ( .IN(n175), .OUT(n176) );
  INVX1 U180 ( .IN(DP_OP_1074_157_5430_n9), .OUT(n177) );
  INVX4 U181 ( .IN(n177), .OUT(n178) );
  NAND2X1 U182 ( .IN1(C2_Z_0), .IN2(DP_OP_1074_157_5430_n33), .OUT(
        DP_OP_1074_157_5430_n31) );
  NAND2X1 U183 ( .IN1(n602), .IN2(n612), .OUT(n248) );
  INVX4 U184 ( .IN(n264), .OUT(n179) );
  NANDX2 U185 ( .IN1(n624), .IN2(C493_DATA2_7), .OUT(n555) );
  NAND2X1 U186 ( .IN1(n624), .IN2(C493_DATA2_4), .OUT(n543) );
  BUF4X U187 ( .IN(DP_OP_1074_157_5430_n10), .OUT(n189) );
  NAND2X1 U188 ( .IN1(n624), .IN2(C493_DATA2_3), .OUT(n625) );
  NAND2X1 U189 ( .IN1(n624), .IN2(C493_DATA2_2), .OUT(n540) );
  BUF4X U190 ( .IN(DP_OP_1074_157_5430_n12), .OUT(n188) );
  NAND2X1 U191 ( .IN1(n624), .IN2(C493_DATA2_1), .OUT(n537) );
  BUF4X U192 ( .IN(DP_OP_1074_157_5430_n13), .OUT(n187) );
  INVX1 U193 ( .IN(n471), .OUT(n128) );
  NANDX2 U194 ( .IN1(n262), .IN2(n1107), .OUT(n468) );
  INVX1 U195 ( .IN(n1114), .OUT(n119) );
  NAND2X1 U196 ( .IN1(n624), .IN2(C493_DATA2_0), .OUT(n552) );
  INVX1 U197 ( .IN(n685), .OUT(n118) );
  NAND2X1 U198 ( .IN1(RSTn), .IN2(n749), .OUT(n410) );
  NAND2X1 U199 ( .IN1(n445), .IN2(n727), .OUT(n367) );
  INVX1 U200 ( .IN(n1110), .OUT(n120) );
  INVX1 U201 ( .IN(n315), .OUT(n316) );
  NANDX2 U202 ( .IN1(n611), .IN2(n628), .OUT(n307) );
  INVX1 U203 ( .IN(n726), .OUT(n634) );
  NAND2X1 U204 ( .IN1(n978), .IN2(n977), .OUT(n1141) );
  INVX4 U205 ( .IN(n309), .OUT(n697) );
  NAND2X1 U206 ( .IN1(n413), .IN2(n412), .OUT(n414) );
  INVX1 U207 ( .IN(n1053), .OUT(n1135) );
  NAND2X1 U208 ( .IN1(n1042), .IN2(n1041), .OUT(n1137) );
  INVX1 U209 ( .IN(n611), .OUT(n630) );
  INVX1 U210 ( .IN(n503), .OUT(n424) );
  INVX1 U211 ( .IN(n1047), .OUT(n1072) );
  NAND2X1 U212 ( .IN1(n745), .IN2(n1067), .OUT(n1019) );
  INVX1 U213 ( .IN(n646), .OUT(n573) );
  NAND2X1 U214 ( .IN1(n386), .IN2(n693), .OUT(n515) );
  NANDX2 U215 ( .IN1(n526), .IN2(n598), .OUT(n312) );
  INVX1 U216 ( .IN(n695), .OUT(n700) );
  INVX1 U217 ( .IN(n453), .OUT(n454) );
  INVX1 U218 ( .IN(n561), .OUT(n638) );
  NAND2X1 U219 ( .IN1(n746), .IN2(n943), .OUT(n1014) );
  INVX1 U220 ( .IN(n1002), .OUT(n1003) );
  INVX1 U221 ( .IN(n357), .OUT(n350) );
  INVX1 U222 ( .IN(n644), .OUT(n567) );
  INVX1 U223 ( .IN(n874), .OUT(n875) );
  INVX1 U224 ( .IN(n668), .OUT(n670) );
  NAND2X1 U225 ( .IN1(n745), .IN2(n1009), .OUT(n1002) );
  INVX1 U226 ( .IN(n678), .OUT(n464) );
  INVX1 U227 ( .IN(n1036), .OUT(n1037) );
  INVX1 U228 ( .IN(n1030), .OUT(n1031) );
  INVX1 U229 ( .IN(n587), .OUT(n641) );
  INVX1 U230 ( .IN(n1018), .OUT(n1022) );
  NAND2X1 U231 ( .IN1(n501), .IN2(n500), .OUT(n502) );
  NAND2X1 U232 ( .IN1(n478), .IN2(n477), .OUT(n479) );
  NANDX2 U233 ( .IN1(n261), .IN2(n244), .OUT(n293) );
  INVX1 U234 ( .IN(n376), .OUT(n373) );
  INVX1 U235 ( .IN(n834), .OUT(n1165) );
  INVX1 U236 ( .IN(n416), .OUT(n417) );
  NANDX2 U237 ( .IN1(n577), .IN2(n576), .OUT(n651) );
  NAND2X1 U238 ( .IN1(n510), .IN2(n511), .OUT(n376) );
  NANDX2 U239 ( .IN1(n193), .IN2(n278), .OUT(n291) );
  NANDX2 U240 ( .IN1(add_x_35_A_8_), .IN2(n1170), .OUT(n1167) );
  NAND2X1 U241 ( .IN1(n261), .IN2(n484), .OUT(n416) );
  INVX4 U242 ( .IN(n1115), .OUT(n755) );
  NANDX2 U243 ( .IN1(n205), .IN2(n639), .OUT(n577) );
  NAND2X1 U244 ( .IN1(n652), .IN2(n1115), .OUT(n579) );
  INVX1 U245 ( .IN(n1068), .OUT(n1069) );
  INVX1 U246 ( .IN(n533), .OUT(n534) );
  NAND2X1 U247 ( .IN1(n257), .IN2(n982), .OUT(n983) );
  INVX4 U248 ( .IN(n1097), .OUT(n712) );
  NANDX2 U249 ( .IN1(n565), .IN2(n564), .OUT(n674) );
  NAND2X1 U250 ( .IN1(n997), .IN2(n982), .OUT(n783) );
  INVX1 U251 ( .IN(n858), .OUT(n1153) );
  NAND2X1 U252 ( .IN1(n1108), .IN2(n791), .OUT(n792) );
  INVX1 U253 ( .IN(n667), .OUT(n744) );
  NAND2X1 U254 ( .IN1(n260), .IN2(n371), .OUT(n418) );
  NANDX2 U255 ( .IN1(carry_reg), .IN2(n268), .OUT(n1097) );
  NANDX2 U256 ( .IN1(n563), .IN2(n562), .OUT(n565) );
  NANDX2 U257 ( .IN1(n202), .IN2(n562), .OUT(n564) );
  NANDX2 U258 ( .IN1(n286), .IN2(n288), .OUT(n331) );
  INVX1 U259 ( .IN(n679), .OUT(n680) );
  NAND2X1 U260 ( .IN1(n808), .IN2(n831), .OUT(n809) );
  NANDX2 U261 ( .IN1(n249), .IN2(n271), .OUT(n699) );
  INVX1 U262 ( .IN(n735), .OUT(ExcCheck_Datain_1_) );
  INVX1 U263 ( .IN(n737), .OUT(ExcCheck_Datain_3_) );
  INVX1 U264 ( .IN(n738), .OUT(ExcCheck_Datain_4_) );
  INVX1 U265 ( .IN(n736), .OUT(ExcCheck_Datain_2_) );
  INVX1 U266 ( .IN(n485), .OUT(n371) );
  INVX1 U267 ( .IN(n740), .OUT(ExcCheck_Datain_6_) );
  NAND2X1 U268 ( .IN1(n1056), .IN2(n1055), .OUT(n1059) );
  INVX1 U269 ( .IN(n739), .OUT(ExcCheck_Datain_5_) );
  INVX1 U270 ( .IN(n794), .OUT(n790) );
  INVX1 U271 ( .IN(n734), .OUT(ExcCheck_Datain_0_) );
  INVX1 U272 ( .IN(n1092), .OUT(n528) );
  INVX1 U273 ( .IN(n531), .OUT(n666) );
  INVX4 U274 ( .IN(n270), .OUT(n271) );
  NAND2X1 U275 ( .IN1(n263), .IN2(n174), .OUT(n282) );
  NANDX2 U276 ( .IN1(n707), .IN2(n269), .OUT(n701) );
  INVX1 U277 ( .IN(n1106), .OUT(n1080) );
  NAND2X1 U278 ( .IN1(n1090), .IN2(n1077), .OUT(n857) );
  NANDX2 U279 ( .IN1(add_x_35_A_4_), .IN2(n1182), .OUT(n1179) );
  INVX1 U280 ( .IN(n253), .OUT(n808) );
  INVX1 U281 ( .IN(n1090), .OUT(n1190) );
  INVX1 U282 ( .IN(n1096), .OUT(n465) );
  NANDX2 U283 ( .IN1(n253), .IN2(Exc_Ack), .OUT(n794) );
  NAND2X1 U284 ( .IN1(n363), .IN2(n1081), .OUT(n448) );
  INVX1 U285 ( .IN(n829), .OUT(n830) );
  INVX1 U286 ( .IN(n815), .OUT(Debug[0]) );
  INVX1 U287 ( .IN(n816), .OUT(Debug[1]) );
  INVX1 U288 ( .IN(n820), .OUT(Debug[4]) );
  INVX1 U289 ( .IN(n817), .OUT(Debug[2]) );
  INVX1 U290 ( .IN(n360), .OUT(n361) );
  INVX1 U291 ( .IN(n370), .OUT(n372) );
  INVX1 U292 ( .IN(n1077), .OUT(n273) );
  NAND2X1 U293 ( .IN1(n836), .IN2(Data_valid), .OUT(n842) );
  NANDX2 U294 ( .IN1(Final_Mantissa_reg[10]), .IN2(n707), .OUT(n270) );
  INVX1 U295 ( .IN(n912), .OUT(n915) );
  INVX4 U296 ( .IN(n760), .OUT(n767) );
  NAND2X1 U297 ( .IN1(n1054), .IN2(n807), .OUT(n831) );
  INVX1 U298 ( .IN(n606), .OUT(n659) );
  INVX1 U299 ( .IN(n818), .OUT(Debug[3]) );
  INVX1 U300 ( .IN(n1100), .OUT(n832) );
  NAND2X1 U301 ( .IN1(RSTn), .IN2(n1100), .OUT(n1077) );
  NANDX2 U302 ( .IN1(n223), .IN2(n1078), .OUT(n1076) );
  NAND2X1 U303 ( .IN1(n259), .IN2(n258), .OUT(n360) );
  INVX1 U304 ( .IN(n1078), .OUT(n272) );
  NANDX2 U305 ( .IN1(add_x_35_A_2_), .IN2(n1118), .OUT(n1185) );
  INVX1 U306 ( .IN(n348), .OUT(n339) );
  NANDX2 U307 ( .IN1(StateMC[2]), .IN2(n845), .OUT(Dataout_valid_BAR) );
  NANDX2 U308 ( .IN1(Datain1[7]), .IN2(n936), .OUT(n774) );
  INVX4 U309 ( .IN(Datain2[7]), .OUT(n936) );
  NANDX2 U310 ( .IN1(StateMC[1]), .IN2(n198), .OUT(n1100) );
  BUF4X U311 ( .IN(Final_Exponent_reg[3]), .OUT(n183) );
  BUF4X U312 ( .IN(Final_Exponent_reg[5]), .OUT(n182) );
  BUF4X U313 ( .IN(Final_Exponent_reg[6]), .OUT(n180) );
  INVX1 U314 ( .IN(n196), .OUT(n186) );
  BUF4X U315 ( .IN(Final_Exponent_reg[0]), .OUT(n181) );
  INVX1 U316 ( .IN(n230), .OUT(n185) );
  INVX4 U317 ( .IN(n205), .OUT(n184) );
  INVX1 U318 ( .IN(n997), .OUT(n984) );
  NAND2X1 U319 ( .IN1(n249), .IN2(n1185), .OUT(n1189) );
  NAND2X1 U320 ( .IN1(n249), .IN2(n1179), .OUT(n1181) );
  NAND2X1 U321 ( .IN1(n249), .IN2(n1173), .OUT(n1175) );
  NAND2X1 U322 ( .IN1(n249), .IN2(n1167), .OUT(n1169) );
  INVX1 U323 ( .IN(n1049), .OUT(n770) );
  NAND2X1 U324 ( .IN1(n1052), .IN2(n940), .OUT(n941) );
  NAND2X1 U325 ( .IN1(n757), .IN2(n1115), .OUT(n1085) );
  INVX1 U326 ( .IN(n432), .OUT(n441) );
  NAND2X1 U327 ( .IN1(n768), .IN2(n774), .OUT(n902) );
  INVX1 U328 ( .IN(n782), .OUT(n781) );
  NAND2X1 U329 ( .IN1(n889), .IN2(n891), .OUT(n890) );
  NAND2X1 U330 ( .IN1(RSTn), .IN2(n1081), .OUT(n1096) );
  NAND2X1 U331 ( .IN1(n802), .IN2(n801), .OUT(n803) );
  INVX1 U332 ( .IN(n648), .OUT(n649) );
  NAND2X1 U333 ( .IN1(n1191), .IN2(n755), .OUT(n730) );
  NANDX2 U334 ( .IN1(n324), .IN2(n636), .OUT(n325) );
  INVX4 U335 ( .IN(n323), .OUT(n324) );
  NANDX2 U336 ( .IN1(n330), .IN2(n636), .OUT(n337) );
  INVX4 U337 ( .IN(n329), .OUT(n330) );
  INVX1 U338 ( .IN(n615), .OUT(n616) );
  NANDX2 U339 ( .IN1(n196), .IN2(n654), .OUT(n656) );
  NAND2X1 U340 ( .IN1(n1115), .IN2(n573), .OUT(n246) );
  INVX4 U341 ( .IN(n1112), .OUT(n733) );
  NANDX2 U342 ( .IN1(n221), .IN2(n268), .OUT(n1112) );
  INVX4 U343 ( .IN(n893), .OUT(n784) );
  NANDX2 U344 ( .IN1(n249), .IN2(n254), .OUT(n1119) );
  NANDX2 U345 ( .IN1(n357), .IN2(n356), .OUT(n693) );
  NANDX2 U346 ( .IN1(n699), .IN2(n666), .OUT(n682) );
  INVX4 U347 ( .IN(n732), .OUT(n355) );
  NAND2X1 U348 ( .IN1(n293), .IN2(n294), .OUT(n311) );
  NAND2X1 U349 ( .IN1(n222), .IN2(n193), .OUT(n243) );
  BUF4X U350 ( .IN(N696), .OUT(n262) );
  NANDX2 U351 ( .IN1(n469), .IN2(n468), .OUT(n470) );
  NANDX2 U352 ( .IN1(n467), .IN2(n466), .OUT(n1123) );
  INVX4 U353 ( .IN(n321), .OUT(n686) );
  NAND2X1 U354 ( .IN1(n262), .IN2(n349), .OUT(n357) );
  INVX4 U355 ( .IN(n1071), .OUT(n745) );
  BUF4X U356 ( .IN(n1186), .OUT(n249) );
  BUF4X U357 ( .IN(n877), .OUT(n255) );
  BUF4X U358 ( .IN(N366), .OUT(n264) );
  INVX4 U359 ( .IN(n498), .OUT(n512) );
  NAND2X1 U360 ( .IN1(n301), .IN2(n525), .OUT(n611) );
  INVX1 U361 ( .IN(n311), .OUT(n526) );
  INVX4 U362 ( .IN(n298), .OUT(n299) );
  NANDX2 U363 ( .IN1(n219), .IN2(n280), .OUT(n298) );
  INVX4 U364 ( .IN(n281), .OUT(n280) );
  INVX4 U365 ( .IN(n1073), .OUT(n746) );
  BUF4X U366 ( .IN(n1187), .OUT(n254) );
  NANDX2 U367 ( .IN1(n379), .IN2(n378), .OUT(n380) );
  BUF4X U368 ( .IN(N152), .OUT(n251) );
  BUF4X U369 ( .IN(N148), .OUT(n252) );
  NANDX2 U370 ( .IN1(n668), .IN2(n743), .OUT(n661) );
  INVX4 U371 ( .IN(n411), .OUT(n386) );
  NANDX2 U372 ( .IN1(n757), .IN2(n730), .OUT(n411) );
  NANDX2 U373 ( .IN1(n757), .IN2(n387), .OUT(n509) );
  INVX4 U374 ( .IN(n1076), .OUT(n757) );
  INVX4 U375 ( .IN(n605), .OUT(C1_Z_1) );
  INVX4 U376 ( .IN(n593), .OUT(C1_Z_2) );
  NAND2X1 U377 ( .IN1(n686), .IN2(n322), .OUT(n725) );
  NANDX2 U378 ( .IN1(n733), .IN2(n637), .OUT(n245) );
  INVX4 U379 ( .IN(n317), .OUT(n318) );
  INVX4 U380 ( .IN(n728), .OUT(n710) );
  NANDX2 U381 ( .IN1(Final_Mantissa_reg[10]), .IN2(n523), .OUT(n295) );
  NANDX2 U382 ( .IN1(n690), .IN2(n331), .OUT(n332) );
  NAND2X1 U383 ( .IN1(n258), .IN2(n285), .OUT(n286) );
  BUF4X U384 ( .IN(n748), .OUT(n250) );
  INVX4 U385 ( .IN(n256), .OUT(n1015) );
  INVX4 U386 ( .IN(n980), .OUT(n1016) );
  NANDX2 U387 ( .IN1(n179), .IN2(n902), .OUT(n980) );
  INVX4 U388 ( .IN(n682), .OUT(n1116) );
  INVX1 U389 ( .IN(n629), .OUT(n658) );
  INVX1 U390 ( .IN(n359), .OUT(n688) );
  NANDX2 U391 ( .IN1(n495), .IN2(n722), .OUT(n352) );
  INVX4 U392 ( .IN(n1108), .OUT(n1088) );
  NANDX2 U393 ( .IN1(n753), .IN2(n757), .OUT(n1104) );
  NAND2X1 U394 ( .IN1(n733), .IN2(n705), .OUT(n696) );
  NANDX2 U395 ( .IN1(n624), .IN2(C493_DATA2_5), .OUT(n546) );
  INVX4 U396 ( .IN(n312), .OUT(n314) );
  INVX4 U397 ( .IN(n434), .OUT(n343) );
  NANDX2 U398 ( .IN1(n259), .IN2(n347), .OUT(n648) );
  INVX4 U399 ( .IN(n572), .OUT(n637) );
  INVX4 U400 ( .IN(n319), .OUT(n320) );
  NANDX2 U401 ( .IN1(n318), .IN2(n331), .OUT(n319) );
  INVX4 U402 ( .IN(n571), .OUT(n574) );
  INVX4 U403 ( .IN(n287), .OUT(n306) );
  NANDX2 U404 ( .IN1(n302), .IN2(n457), .OUT(n446) );
  NANDX2 U405 ( .IN1(n195), .IN2(n279), .OUT(n281) );
  INVX4 U406 ( .IN(n294), .OUT(n279) );
  INVX4 U407 ( .IN(n295), .OUT(n296) );
  NANDX2 U408 ( .IN1(n204), .IN2(n292), .OUT(n294) );
  INVX4 U409 ( .IN(n243), .OUT(n242) );
  NANDX2 U410 ( .IN1(n203), .IN2(n276), .OUT(n289) );
  INVX4 U411 ( .IN(n288), .OUT(n276) );
  INVX4 U412 ( .IN(n332), .OUT(n333) );
  INVX4 U413 ( .IN(n285), .OUT(n275) );
  NANDX2 U414 ( .IN1(n190), .IN2(n362), .OUT(n285) );
  NANDX2 U415 ( .IN1(n559), .IN2(n558), .OUT(n560) );
  NANDX2 U416 ( .IN1(n755), .IN2(n534), .OUT(n535) );
  NAND2X1 U417 ( .IN1(carry_reg), .IN2(n1095), .OUT(n466) );
  INVX4 U418 ( .IN(n742), .OUT(ExcCheck_Datain_14_) );
  INVX4 U419 ( .IN(n741), .OUT(ExcCheck_Datain_12_) );
  INVX4 U420 ( .IN(n822), .OUT(ExcCheck_Datain_11_) );
  INVX4 U421 ( .IN(n827), .OUT(ExcCheck_Datain_9_) );
  INVX4 U422 ( .IN(n824), .OUT(ExcCheck_Datain_8_) );
  NAND2X1 U423 ( .IN1(n198), .IN2(n223), .OUT(n860) );
  NANDX2 U424 ( .IN1(n1034), .IN2(n1033), .OUT(n1138) );
  NANDX2 U425 ( .IN1(n1064), .IN2(n1063), .OUT(n1134) );
  INVX4 U426 ( .IN(n1050), .OUT(n1061) );
  INVX4 U427 ( .IN(n1119), .OUT(n1070) );
  INVX4 U428 ( .IN(n850), .OUT(n856) );
  INVX1 U429 ( .IN(Mode[1]), .OUT(n814) );
  INVX4 U430 ( .IN(n804), .OUT(n825) );
  NANDX2 U431 ( .IN1(n973), .IN2(n980), .OUT(n1039) );
  NANDX2 U432 ( .IN1(n952), .IN2(n951), .OUT(n966) );
  NANDX2 U433 ( .IN1(n969), .IN2(n968), .OUT(n1007) );
  INVX4 U434 ( .IN(n257), .OUT(n979) );
  INVX4 U435 ( .IN(n415), .OUT(n406) );
  INVX4 U436 ( .IN(n426), .OUT(n409) );
  NAND2X1 U437 ( .IN1(Datain1[7]), .IN2(n745), .OUT(n553) );
  NANDX2 U438 ( .IN1(n395), .IN2(n394), .OUT(n396) );
  NANDX2 U439 ( .IN1(n369), .IN2(n368), .OUT(n442) );
  INVX4 U440 ( .IN(n433), .OUT(n439) );
  NANDX2 U441 ( .IN1(n384), .IN2(n383), .OUT(n433) );
  NANDX2 U442 ( .IN1(n428), .IN2(n427), .OUT(n429) );
  NANDX2 U443 ( .IN1(n402), .IN2(n401), .OUT(n415) );
  NANDX2 U444 ( .IN1(n400), .IN2(n399), .OUT(n426) );
  INVX4 U445 ( .IN(n251), .OUT(N168) );
  NANDX2 U446 ( .IN1(n251), .IN2(n1067), .OUT(n1047) );
  INVX4 U447 ( .IN(n949), .OUT(n1001) );
  NANDX2 U448 ( .IN1(N156), .IN2(n1040), .OUT(n949) );
  INVX4 U449 ( .IN(n950), .OUT(n1040) );
  NANDX2 U450 ( .IN1(n1075), .IN2(n947), .OUT(n950) );
  INVX4 U451 ( .IN(n1065), .OUT(n1075) );
  INVX4 U452 ( .IN(n929), .OUT(n992) );
  INVX4 U453 ( .IN(n909), .OUT(n927) );
  BUF4X U454 ( .IN(Datain1[6]), .OUT(n257) );
  BUF4X U455 ( .IN(Datain1[5]), .OUT(n256) );
  NANDX2 U456 ( .IN1(n767), .IN2(n774), .OUT(N366) );
  NANDX2 U457 ( .IN1(n997), .IN2(n946), .OUT(n1065) );
  NANDX2 U458 ( .IN1(n888), .IN2(n919), .OUT(n891) );
  INVX4 U459 ( .IN(n777), .OUT(n776) );
  INVX4 U460 ( .IN(n1051), .OUT(n1028) );
  NANDX2 U461 ( .IN1(n747), .IN2(n1193), .OUT(n1051) );
  INVX4 U462 ( .IN(n514), .OUT(n504) );
  NANDX2 U463 ( .IN1(n1096), .IN2(n1092), .OUT(n679) );
  NANDX2 U464 ( .IN1(n671), .IN2(n800), .OUT(n673) );
  NANDX2 U465 ( .IN1(n650), .IN2(n649), .OUT(n668) );
  NANDX2 U466 ( .IN1(n263), .IN2(n463), .OUT(n678) );
  INVX4 U467 ( .IN(n455), .OUT(n364) );
  INVX4 U468 ( .IN(n410), .OUT(n527) );
  INVX4 U469 ( .IN(n482), .OUT(n749) );
  NANDX2 U470 ( .IN1(n493), .IN2(n491), .OUT(n482) );
  NANDX2 U471 ( .IN1(n273), .IN2(n272), .OUT(n1092) );
  NANDX2 U472 ( .IN1(n337), .IN2(n491), .OUT(n336) );
  NANDX2 U473 ( .IN1(n733), .IN2(n757), .OUT(n1099) );
  NANDX2 U474 ( .IN1(n1083), .IN2(n1082), .OUT(n1084) );
  INVX4 U475 ( .IN(n366), .OUT(n689) );
  NANDX2 U476 ( .IN1(n354), .IN2(n353), .OUT(n520) );
  INVX4 U477 ( .IN(n476), .OUT(n750) );
  INVX4 U478 ( .IN(n519), .OUT(n487) );
  INVX4 U479 ( .IN(n382), .OUT(n521) );
  NANDX2 U480 ( .IN1(n386), .IN2(n695), .OUT(n382) );
  INVX4 U481 ( .IN(n488), .OUT(n754) );
  INVX4 U482 ( .IN(n352), .OUT(n518) );
  NANDX2 U483 ( .IN1(n681), .IN2(n722), .OUT(n519) );
  INVX4 U484 ( .IN(n1104), .OUT(n513) );
  NANDX2 U485 ( .IN1(n497), .IN2(n496), .OUT(n514) );
  INVX1 U486 ( .IN(Adder_ack), .OUT(n807) );
  INVX4 U487 ( .IN(n448), .OUT(n511) );
  NANDX2 U488 ( .IN1(n372), .IN2(n484), .OUT(n510) );
  INVX4 U489 ( .IN(n418), .OUT(n484) );
  NANDX2 U490 ( .IN1(n495), .IN2(n496), .OUT(n476) );
  INVX4 U491 ( .IN(n722), .OUT(n496) );
  NANDX2 U492 ( .IN1(n351), .IN2(n646), .OUT(n722) );
  INVX4 U493 ( .IN(n681), .OUT(n495) );
  NANDX2 U494 ( .IN1(n358), .IN2(n1086), .OUT(n488) );
  INVX4 U495 ( .IN(n693), .OUT(n1086) );
  NANDX2 U496 ( .IN1(n713), .IN2(n355), .OUT(n695) );
  NANDX2 U497 ( .IN1(n587), .IN2(n648), .OUT(n732) );
  NANDX2 U498 ( .IN1(n493), .IN2(n492), .OUT(n508) );
  INVX4 U499 ( .IN(n328), .OUT(n492) );
  NANDX2 U500 ( .IN1(n752), .IN2(n727), .OUT(n473) );
  NANDX2 U501 ( .IN1(n365), .IN2(n752), .OUT(n327) );
  NANDX2 U502 ( .IN1(n572), .IN2(n326), .OUT(n445) );
  INVX4 U503 ( .IN(n325), .OUT(n326) );
  NANDX2 U504 ( .IN1(n717), .IN2(n316), .OUT(n365) );
  INVX4 U505 ( .IN(n307), .OUT(n717) );
  INVX4 U506 ( .IN(n337), .OUT(n493) );
  NAND2X1 U507 ( .IN1(Datain1[8]), .IN2(n745), .OUT(n538) );
  NAND2X1 U508 ( .IN1(Datain1[9]), .IN2(n745), .OUT(n541) );
  NAND2X1 U509 ( .IN1(Datain1[10]), .IN2(n745), .OUT(n626) );
  NAND2X1 U510 ( .IN1(Datain1[11]), .IN2(n745), .OUT(n544) );
  NANDX2 U511 ( .IN1(n624), .IN2(C493_DATA2_6), .OUT(n549) );
  NAND2X1 U512 ( .IN1(Datain1[13]), .IN2(n745), .OUT(n550) );
  INVX4 U513 ( .IN(n607), .OUT(n609) );
  NANDX2 U514 ( .IN1(n659), .IN2(n629), .OUT(n607) );
  NANDX2 U515 ( .IN1(n247), .IN2(n601), .OUT(n603) );
  INVX4 U516 ( .IN(n248), .OUT(n247) );
  NANDX2 U517 ( .IN1(n314), .IN2(n313), .OUT(n632) );
  NANDX2 U518 ( .IN1(n594), .IN2(n656), .OUT(n660) );
  INVX4 U519 ( .IN(n656), .OUT(n631) );
  NANDX2 U520 ( .IN1(n591), .IN2(n619), .OUT(n604) );
  NANDX2 U521 ( .IN1(n590), .IN2(n589), .OUT(n619) );
  NANDX2 U522 ( .IN1(n343), .IN2(n347), .OUT(n587) );
  NANDX2 U523 ( .IN1(n692), .IN2(n334), .OUT(n636) );
  INVX4 U524 ( .IN(n640), .OUT(n590) );
  NANDX2 U525 ( .IN1(n586), .IN2(n635), .OUT(n640) );
  INVX4 U526 ( .IN(n635), .OUT(n650) );
  NANDX2 U527 ( .IN1(n582), .IN2(n639), .OUT(n635) );
  NANDX2 U528 ( .IN1(n633), .IN2(n580), .OUT(n615) );
  NANDX2 U529 ( .IN1(n310), .IN2(n697), .OUT(n708) );
  INVX4 U530 ( .IN(n651), .OUT(n633) );
  NANDX2 U531 ( .IN1(n524), .IN2(n697), .OUT(n726) );
  INVX4 U532 ( .IN(n308), .OUT(n524) );
  INVX4 U533 ( .IN(n577), .OUT(n654) );
  NANDX2 U534 ( .IN1(n574), .IN2(n601), .OUT(C1_Z_3) );
  NANDX2 U535 ( .IN1(n647), .IN2(n675), .OUT(n601) );
  NANDX2 U536 ( .IN1(n246), .IN2(n245), .OUT(n675) );
  NANDX2 U537 ( .IN1(n320), .IN2(n334), .OUT(n572) );
  NANDX2 U538 ( .IN1(n350), .IN2(n356), .OUT(n646) );
  INVX4 U539 ( .IN(n731), .OUT(n356) );
  NANDX2 U540 ( .IN1(n644), .IN2(n561), .OUT(n731) );
  INVX4 U541 ( .IN(n674), .OUT(n647) );
  NANDX2 U542 ( .IN1(n643), .IN2(n569), .OUT(n618) );
  NANDX2 U543 ( .IN1(n346), .IN2(n349), .OUT(n644) );
  NANDX2 U544 ( .IN1(n306), .IN2(n334), .OUT(n628) );
  NANDX2 U545 ( .IN1(n284), .IN2(n283), .OUT(n499) );
  NANDX2 U546 ( .IN1(n566), .IN2(n674), .OUT(n643) );
  NANDX2 U547 ( .IN1(n333), .IN2(n334), .OUT(n728) );
  NANDX2 U548 ( .IN1(n321), .IN2(n322), .OUT(n305) );
  NANDX2 U549 ( .IN1(n303), .IN2(n313), .OUT(n309) );
  INVX4 U550 ( .IN(n446), .OUT(n313) );
  INVX4 U551 ( .IN(n724), .OUT(n457) );
  NANDX2 U552 ( .IN1(n301), .IN2(n300), .OUT(n724) );
  INVX4 U553 ( .IN(n297), .OUT(n303) );
  NANDX2 U554 ( .IN1(n311), .IN2(n598), .OUT(n297) );
  NANDX2 U555 ( .IN1(n296), .IN2(n302), .OUT(n598) );
  INVX4 U556 ( .IN(n244), .OUT(n292) );
  NANDX2 U557 ( .IN1(n242), .IN2(n278), .OUT(n244) );
  NANDX2 U558 ( .IN1(n359), .IN2(n308), .OUT(n304) );
  NANDX2 U559 ( .IN1(n290), .IN2(n291), .OUT(n359) );
  INVX4 U560 ( .IN(n289), .OUT(n278) );
  INVX4 U561 ( .IN(n474), .OUT(n690) );
  NANDX2 U562 ( .IN1(n263), .IN2(n349), .OUT(n561) );
  INVX4 U563 ( .IN(n345), .OUT(n349) );
  NANDX2 U564 ( .IN1(n344), .IN2(n347), .OUT(n345) );
  INVX4 U565 ( .IN(n729), .OUT(n347) );
  NANDX2 U566 ( .IN1(n342), .IN2(n713), .OUT(n729) );
  INVX4 U567 ( .IN(n341), .OUT(n713) );
  NANDX2 U568 ( .IN1(n578), .IN2(n575), .OUT(n341) );
  NANDX2 U569 ( .IN1(n260), .IN2(n342), .OUT(n575) );
  NANDX2 U570 ( .IN1(n340), .IN2(n342), .OUT(n578) );
  INVX4 U571 ( .IN(n698), .OUT(n342) );
  NANDX2 U572 ( .IN1(n714), .IN2(n339), .OUT(n698) );
  INVX4 U573 ( .IN(n338), .OUT(n714) );
  BUF4X U574 ( .IN(Final_Mantissa_reg[3]), .OUT(n258) );
  BUF4X U575 ( .IN(Final_Mantissa_reg[4]), .OUT(n259) );
  INVX4 U576 ( .IN(n564), .OUT(n639) );
  INVX4 U577 ( .IN(n560), .OUT(n562) );
  NANDX2 U578 ( .IN1(n535), .IN2(n250), .OUT(n536) );
  NANDX2 U579 ( .IN1(n532), .IN2(n531), .OUT(n667) );
  NANDX2 U580 ( .IN1(n756), .IN2(n271), .OUT(n1191) );
  INVX4 U581 ( .IN(n249), .OUT(n756) );
  NANDX2 U582 ( .IN1(n701), .IN2(n1097), .OUT(n1115) );
  INVX4 U583 ( .IN(n267), .OUT(n268) );
  NANDX2 U584 ( .IN1(n249), .IN2(n270), .OUT(n267) );
  NAND2X1 U585 ( .IN1(Datain1[14]), .IN2(n745), .OUT(n556) );
  NANDX2 U586 ( .IN1(n843), .IN2(n844), .OUT(n1071) );
  INVX1 U587 ( .IN(Datain1[14]), .OUT(n885) );
  NAND2X1 U588 ( .IN1(Datain1[14]), .IN2(n886), .OUT(n841) );
  INVX1 U589 ( .IN(Datain2[14]), .OUT(n886) );
  INVX1 U590 ( .IN(Datain2[13]), .OUT(n840) );
  INVX1 U591 ( .IN(Datain2[12]), .OUT(n932) );
  INVX1 U592 ( .IN(Datain1[11]), .OUT(n892) );
  NAND2X1 U593 ( .IN1(Datain1[8]), .IN2(n935), .OUT(n775) );
  INVX1 U594 ( .IN(Datain2[8]), .OUT(n935) );
  INVX1 U595 ( .IN(Datain1[9]), .OUT(n870) );
  INVX1 U596 ( .IN(Datain2[9]), .OUT(n763) );
  INVX1 U597 ( .IN(Datain2[11]), .OUT(n933) );
  NANDX2 U598 ( .IN1(n530), .IN2(n747), .OUT(n623) );
  NAND2X1 U599 ( .IN1(RSTn), .IN2(n836), .OUT(n837) );
  NAND2X1 U600 ( .IN1(n223), .IN2(n199), .OUT(n838) );
  INVX4 U601 ( .IN(RSTn), .OUT(n265) );
  NAND2X1 U602 ( .IN1(n733), .IN2(n697), .OUT(n706) );
  INVX1 U603 ( .IN(n719), .OUT(n720) );
  INVX1 U604 ( .IN(n707), .OUT(n721) );
  NAND2X1 U605 ( .IN1(n1088), .IN2(Adder_dataout[5]), .OUT(n375) );
  INVX1 U606 ( .IN(n489), .OUT(n481) );
  INVX1 U607 ( .IN(n491), .OUT(n506) );
  NAND2X1 U608 ( .IN1(Final_Mantissa_reg[10]), .IN2(Final_Mantissa_reg[9]), 
        .OUT(n447) );
  BUF4X U609 ( .IN(n826), .OUT(n253) );
  NAND2X1 U610 ( .IN1(n445), .IN2(n365), .OUT(n366) );
  NAND2X1 U611 ( .IN1(Adder_ack), .IN2(n1054), .OUT(n1108) );
  NAND2X1 U612 ( .IN1(Final_Mantissa_reg[5]), .IN2(n361), .OUT(n485) );
  NAND2X1 U613 ( .IN1(Final_Mantissa_reg[8]), .IN2(n261), .OUT(n370) );
  INVX1 U614 ( .IN(n696), .OUT(n387) );
  NAND2X1 U615 ( .IN1(Datain1[12]), .IN2(n745), .OUT(n547) );
  INVX1 U616 ( .IN(n302), .OUT(n525) );
  NAND2X1 U617 ( .IN1(n220), .IN2(n631), .OUT(n629) );
  NAND2X1 U618 ( .IN1(Final_Mantissa_reg[9]), .IN2(n194), .OUT(n606) );
  INVX1 U619 ( .IN(n701), .OUT(n610) );
  NAND2X1 U620 ( .IN1(n220), .IN2(n654), .OUT(n594) );
  INVX1 U621 ( .IN(n598), .OUT(n723) );
  NAND2X1 U622 ( .IN1(Final_Mantissa_reg[8]), .IN2(n714), .OUT(n655) );
  NAND2X1 U623 ( .IN1(n1115), .IN2(n641), .OUT(n588) );
  NAND2X1 U624 ( .IN1(n258), .IN2(n203), .OUT(n434) );
  NAND2X1 U625 ( .IN1(n220), .IN2(n639), .OUT(n586) );
  INVX1 U626 ( .IN(n725), .OUT(n583) );
  NAND2X1 U627 ( .IN1(Final_Exponent_reg[1]), .IN2(n184), .OUT(n582) );
  INVX1 U628 ( .IN(n578), .OUT(n652) );
  INVX1 U629 ( .IN(n575), .OUT(n653) );
  NAND2X1 U630 ( .IN1(n1115), .IN2(n567), .OUT(n568) );
  NAND2X1 U631 ( .IN1(n262), .IN2(n192), .OUT(n283) );
  NAND2X1 U632 ( .IN1(Final_Mantissa_reg[1]), .IN2(n197), .OUT(n284) );
  NAND2X1 U633 ( .IN1(n181), .IN2(n183), .OUT(n566) );
  NAND2X1 U634 ( .IN1(Final_Mantissa_reg[5]), .IN2(n289), .OUT(n290) );
  NAND2X1 U635 ( .IN1(n285), .IN2(n282), .OUT(n474) );
  NAND2X1 U636 ( .IN1(n195), .IN2(n204), .OUT(n348) );
  NAND2X1 U637 ( .IN1(n194), .IN2(n219), .OUT(n338) );
  INVX1 U638 ( .IN(n844), .OUT(n529) );
  NAND2X1 U639 ( .IN1(carry_reg), .IN2(n206), .OUT(n266) );
  BUF4X U640 ( .IN(Final_Mantissa_reg[2]), .OUT(n263) );
  BUF4X U641 ( .IN(Final_Mantissa_reg[7]), .OUT(n261) );
  BUF4X U642 ( .IN(Final_Mantissa_reg[6]), .OUT(n260) );
  MUX2X1 U643 ( .IN1(Final_Mantissa_reg[8]), .IN2(n195), .S(n294), .OUT(n523)
         );
  TIEHI U644 ( .OUT(n73) );
  NAND2X1 U645 ( .IN1(n513), .IN2(n523), .OUT(n378) );
  INVX4 U646 ( .IN(n252), .OUT(N156) );
  INVX4 U647 ( .IN(n254), .OUT(n1091) );
  MUX2X1 U648 ( .IN1(n191), .IN2(n216), .S(n215), .OUT(n1186) );
  OAI21 U649 ( .IN1(carry_reg), .IN2(n206), .IN3(n266), .OUT(n707) );
  NOR2X1 U650 ( .IN1(Final_Mantissa_reg[10]), .IN2(n249), .OUT(n269) );
  INVX4 U651 ( .IN(n699), .OUT(n753) );
  NANDX2 U652 ( .IN1(n201), .IN2(n275), .OUT(n288) );
  MUX2X1 U653 ( .IN1(n219), .IN2(Final_Mantissa_reg[9]), .S(n281), .OUT(n302)
         );
  NAND3X1 U654 ( .IN1(n474), .IN2(n499), .IN3(n331), .OUT(n287) );
  MUX2X1 U655 ( .IN1(n203), .IN2(n259), .S(n288), .OUT(n321) );
  MUX2X1 U656 ( .IN1(n222), .IN2(n260), .S(n291), .OUT(n308) );
  NOR2X1 U657 ( .IN1(n304), .IN2(n309), .OUT(n322) );
  INVX4 U658 ( .IN(n305), .OUT(n334) );
  NOR2X1 U659 ( .IN1(n359), .IN2(n524), .OUT(n310) );
  INVX4 U660 ( .IN(n331), .OUT(n692) );
  NAND3X1 U661 ( .IN1(n708), .IN2(n632), .IN3(n636), .OUT(n315) );
  NAND3X1 U662 ( .IN1(n262), .IN2(n263), .IN3(Final_Mantissa_reg[1]), .OUT(
        n317) );
  NAND3X1 U663 ( .IN1(n173), .IN2(n632), .IN3(n725), .OUT(n323) );
  INVX4 U664 ( .IN(n445), .OUT(n752) );
  INVX4 U665 ( .IN(n327), .OUT(n687) );
  INVX4 U666 ( .IN(n365), .OUT(n727) );
  INVX4 U667 ( .IN(n473), .OUT(n751) );
  AOI22 U668 ( .IN1(n687), .IN2(n262), .IN3(n499), .IN4(n751), .OUT(n328) );
  NAND3X1 U669 ( .IN1(n708), .IN2(n726), .IN3(n725), .OUT(n329) );
  NAND3X1 U670 ( .IN1(n258), .IN2(n262), .IN3(n334), .OUT(n335) );
  NAND3X1 U671 ( .IN1(n728), .IN2(n628), .IN3(n335), .OUT(n705) );
  NOR2X1 U672 ( .IN1(n1099), .IN2(n705), .OUT(n491) );
  INVX4 U673 ( .IN(n336), .OUT(n522) );
  NOR2X1 U674 ( .IN1(n260), .IN2(n193), .OUT(n340) );
  NOR2X1 U675 ( .IN1(n263), .IN2(n192), .OUT(n346) );
  NOR2X1 U676 ( .IN1(n259), .IN2(n258), .OUT(n344) );
  AOI21 U677 ( .IN1(n714), .IN2(n348), .IN3(n732), .OUT(n351) );
  NOR2X1 U678 ( .IN1(n495), .IN2(n722), .OUT(n517) );
  AOI22 U679 ( .IN1(n518), .IN2(n258), .IN3(n259), .IN4(n517), .OUT(n354) );
  AOI22 U680 ( .IN1(n263), .IN2(n487), .IN3(Final_Mantissa_reg[5]), .IN4(n750), 
        .OUT(n353) );
  NOR2X1 U681 ( .IN1(n411), .IN2(n695), .OUT(n358) );
  NOR2X1 U682 ( .IN1(n249), .IN2(n707), .OUT(n531) );
  NOR2X1 U683 ( .IN1(n666), .IN2(n1076), .OUT(n498) );
  AOI21 U684 ( .IN1(n362), .IN2(n201), .IN3(n190), .OUT(n363) );
  OAI21 U685 ( .IN1(n265), .IN2(n364), .IN3(n1092), .OUT(n490) );
  AOI22 U686 ( .IN1(n689), .IN2(n499), .IN3(n692), .IN4(n687), .OUT(n369) );
  INVX4 U687 ( .IN(n367), .OUT(n691) );
  AOI22 U688 ( .IN1(n691), .IN2(n690), .IN3(n751), .IN4(n686), .OUT(n368) );
  NOR2X1 U689 ( .IN1(n373), .IN2(n455), .OUT(n374) );
  OAI21 U690 ( .IN1(n488), .IN2(n476), .IN3(n374), .OUT(n516) );
  OAI21 U691 ( .IN1(n416), .IN2(n376), .IN3(n375), .OUT(n377) );
  AOI21 U692 ( .IN1(n498), .IN2(Final_Mantissa_reg[9]), .IN3(n377), .OUT(n379)
         );
  AOI21 U693 ( .IN1(n516), .IN2(Final_Mantissa_reg[8]), .IN3(n380), .OUT(n392)
         );
  AOI22 U694 ( .IN1(n518), .IN2(n260), .IN3(n261), .IN4(n517), .OUT(n381) );
  OAI21 U695 ( .IN1(n193), .IN2(n519), .IN3(n381), .OUT(n385) );
  AOI22 U696 ( .IN1(n518), .IN2(n263), .IN3(n258), .IN4(n517), .OUT(n384) );
  AOI22 U697 ( .IN1(Final_Mantissa_reg[1]), .IN2(n487), .IN3(n259), .IN4(n750), 
        .OUT(n383) );
  AOI22 U698 ( .IN1(n385), .IN2(n754), .IN3(n521), .IN4(n433), .OUT(n391) );
  NOR2X1 U699 ( .IN1(n515), .IN2(n476), .OUT(n389) );
  NOR2X1 U700 ( .IN1(n509), .IN2(n473), .OUT(n388) );
  OAI21 U701 ( .IN1(n389), .IN2(n388), .IN3(n262), .OUT(n390) );
  NAND3X1 U702 ( .IN1(n392), .IN2(n391), .IN3(n390), .OUT(n393) );
  AOI21 U703 ( .IN1(n442), .IN2(n522), .IN3(n393), .OUT(n398) );
  AOI22 U704 ( .IN1(n689), .IN2(n688), .IN3(n526), .IN4(n687), .OUT(n395) );
  AOI22 U705 ( .IN1(n691), .IN2(n524), .IN3(n751), .IN4(n523), .OUT(n394) );
  AOI22 U706 ( .IN1(Final_Mantissa_reg[8]), .IN2(n528), .IN3(n396), .IN4(n527), 
        .OUT(n397) );
  OAI21 U707 ( .IN1(n265), .IN2(n398), .IN3(n397), .OUT(n1126) );
  AOI22 U708 ( .IN1(n689), .IN2(n262), .IN3(n690), .IN4(n687), .OUT(n400) );
  AOI22 U709 ( .IN1(n691), .IN2(n499), .IN3(n692), .IN4(n751), .OUT(n399) );
  AOI22 U710 ( .IN1(n487), .IN2(n262), .IN3(Final_Mantissa_reg[1]), .IN4(n518), 
        .OUT(n402) );
  AOI22 U711 ( .IN1(n263), .IN2(n517), .IN3(n258), .IN4(n750), .OUT(n401) );
  AOI22 U712 ( .IN1(Adder_dataout[0]), .IN2(n1088), .IN3(n201), .IN4(n511), 
        .OUT(n403) );
  OAI21 U713 ( .IN1(n203), .IN2(n512), .IN3(n403), .OUT(n404) );
  AOI21 U714 ( .IN1(n692), .IN2(n513), .IN3(n404), .OUT(n405) );
  OAI21 U715 ( .IN1(n488), .IN2(n406), .IN3(n405), .OUT(n407) );
  AOI22 U716 ( .IN1(n258), .IN2(n490), .IN3(RSTn), .IN4(n407), .OUT(n408) );
  OAI21 U717 ( .IN1(n410), .IN2(n409), .IN3(n408), .OUT(n1131) );
  NOR2X1 U718 ( .IN1(n411), .IN2(n693), .OUT(n503) );
  AOI22 U719 ( .IN1(n517), .IN2(n260), .IN3(Final_Mantissa_reg[5]), .IN4(n518), 
        .OUT(n413) );
  AOI22 U720 ( .IN1(n259), .IN2(n487), .IN3(n261), .IN4(n750), .OUT(n412) );
  AOI21 U721 ( .IN1(n415), .IN2(n695), .IN3(n414), .OUT(n423) );
  AOI21 U722 ( .IN1(n418), .IN2(n204), .IN3(n417), .OUT(n419) );
  AOI22 U723 ( .IN1(n1088), .IN2(Adder_dataout[4]), .IN3(n511), .IN4(n419), 
        .OUT(n420) );
  OAI21 U724 ( .IN1(n195), .IN2(n512), .IN3(n420), .OUT(n421) );
  AOI21 U725 ( .IN1(n526), .IN2(n513), .IN3(n421), .OUT(n422) );
  OAI21 U726 ( .IN1(n424), .IN2(n423), .IN3(n422), .OUT(n425) );
  AOI21 U727 ( .IN1(n426), .IN2(n522), .IN3(n425), .OUT(n431) );
  AOI22 U728 ( .IN1(n689), .IN2(n686), .IN3(n524), .IN4(n687), .OUT(n428) );
  AOI22 U729 ( .IN1(n691), .IN2(n688), .IN3(n526), .IN4(n751), .OUT(n427) );
  AOI22 U730 ( .IN1(n261), .IN2(n490), .IN3(n429), .IN4(n527), .OUT(n430) );
  OAI21 U731 ( .IN1(n265), .IN2(n431), .IN3(n430), .OUT(n1127) );
  AOI22 U732 ( .IN1(n750), .IN2(n521), .IN3(n751), .IN4(n522), .OUT(n432) );
  OAI21 U733 ( .IN1(n258), .IN2(n203), .IN3(n434), .OUT(n435) );
  AOI22 U734 ( .IN1(n1088), .IN2(Adder_dataout[1]), .IN3(n435), .IN4(n511), 
        .OUT(n436) );
  OAI21 U735 ( .IN1(n193), .IN2(n512), .IN3(n436), .OUT(n437) );
  AOI21 U736 ( .IN1(n513), .IN2(n686), .IN3(n437), .OUT(n438) );
  OAI21 U737 ( .IN1(n488), .IN2(n439), .IN3(n438), .OUT(n440) );
  AOI21 U738 ( .IN1(n441), .IN2(n262), .IN3(n440), .OUT(n444) );
  AOI22 U739 ( .IN1(n259), .IN2(n490), .IN3(n527), .IN4(n442), .OUT(n443) );
  OAI21 U740 ( .IN1(n265), .IN2(n444), .IN3(n443), .OUT(n1130) );
  OAI21 U741 ( .IN1(n446), .IN2(n445), .IN3(n749), .OUT(n460) );
  OAI21 U742 ( .IN1(n219), .IN2(n510), .IN3(n194), .OUT(n450) );
  NOR2X1 U743 ( .IN1(n447), .IN2(n510), .OUT(n463) );
  NOR2X1 U744 ( .IN1(n448), .IN2(n463), .OUT(n449) );
  AOI22 U745 ( .IN1(n1088), .IN2(Adder_dataout[7]), .IN3(n450), .IN4(n449), 
        .OUT(n451) );
  OAI21 U746 ( .IN1(n1076), .IN2(n1191), .IN3(n451), .OUT(n452) );
  AOI21 U747 ( .IN1(carry_reg), .IN2(n498), .IN3(n452), .OUT(n453) );
  AOI21 U748 ( .IN1(Final_Mantissa_reg[10]), .IN2(n455), .IN3(n454), .OUT(n456) );
  OAI21 U749 ( .IN1(n1104), .IN2(n457), .IN3(n456), .OUT(n458) );
  NOR2X1 U750 ( .IN1(n458), .IN2(n522), .OUT(n459) );
  NAND3X1 U751 ( .IN1(n509), .IN2(n460), .IN3(n459), .OUT(n461) );
  OAI21 U752 ( .IN1(n461), .IN2(n1089), .IN3(RSTn), .OUT(n462) );
  OAI21 U753 ( .IN1(n1092), .IN2(n194), .IN3(n462), .OUT(n1124) );
  AOI22 U754 ( .IN1(Adder_carryout), .IN2(n1094), .IN3(n465), .IN4(n464), 
        .OUT(n467) );
  AOI22 U755 ( .IN1(Final_Mantissa_reg[1]), .IN2(n498), .IN3(n200), .IN4(n1088), .OUT(n469) );
  AOI22 U756 ( .IN1(n262), .IN2(n679), .IN3(RSTn), .IN4(n470), .OUT(n471) );
  AOI22 U757 ( .IN1(n687), .IN2(n499), .IN3(n262), .IN4(n691), .OUT(n472) );
  OAI21 U758 ( .IN1(n474), .IN2(n473), .IN3(n472), .OUT(n489) );
  AOI22 U759 ( .IN1(n517), .IN2(Final_Mantissa_reg[1]), .IN3(n262), .IN4(n518), 
        .OUT(n475) );
  OAI21 U760 ( .IN1(n190), .IN2(n476), .IN3(n475), .OUT(n486) );
  AOI22 U761 ( .IN1(n263), .IN2(n1080), .IN3(n258), .IN4(n498), .OUT(n478) );
  AOI22 U762 ( .IN1(n1088), .IN2(n237), .IN3(n690), .IN4(n513), .OUT(n477) );
  AOI21 U763 ( .IN1(n486), .IN2(n754), .IN3(n479), .OUT(n480) );
  OAI21 U764 ( .IN1(n482), .IN2(n481), .IN3(n480), .OUT(n483) );
  AOI22 U765 ( .IN1(n263), .IN2(n679), .IN3(RSTn), .IN4(n483), .OUT(n665) );
  OAI21 U766 ( .IN1(n262), .IN2(n495), .IN3(n700), .OUT(n494) );
  AOI21 U767 ( .IN1(n495), .IN2(n192), .IN3(n494), .OUT(n497) );
  AOI22 U768 ( .IN1(Final_Mantissa_reg[1]), .IN2(n1080), .IN3(n263), .IN4(n498), .OUT(n501) );
  AOI22 U769 ( .IN1(n1088), .IN2(n238), .IN3(n499), .IN4(n513), .OUT(n500) );
  AOI21 U770 ( .IN1(n504), .IN2(n503), .IN3(n502), .OUT(n505) );
  OAI21 U771 ( .IN1(n506), .IN2(n508), .IN3(n505), .OUT(n507) );
  AOI22 U772 ( .IN1(Final_Mantissa_reg[1]), .IN2(n679), .IN3(RSTn), .IN4(n507), 
        .OUT(n672) );
  NOR2X1 U773 ( .IN1(n265), .IN2(n1076), .OUT(n748) );
  INVX4 U774 ( .IN(n250), .OUT(n1193) );
  NANDX2 U775 ( .IN1(n843), .IN2(n529), .OUT(n1073) );
  OAI21 U776 ( .IN1(n753), .IN2(n835), .IN3(n250), .OUT(n530) );
  AOI21 U777 ( .IN1(RSTn), .IN2(n838), .IN3(n859), .OUT(n747) );
  AOI22 U778 ( .IN1(n186), .IN2(n623), .IN3(Datain2[8]), .IN4(n746), .OUT(n539) );
  NAND3X1 U779 ( .IN1(n1191), .IN2(n667), .IN3(n1112), .OUT(n533) );
  INVX4 U780 ( .IN(n536), .OUT(n624) );
  NAND3X1 U781 ( .IN1(n539), .IN2(n538), .IN3(n537), .OUT(n1157) );
  AOI22 U782 ( .IN1(n184), .IN2(n623), .IN3(Datain2[9]), .IN4(n746), .OUT(n542) );
  NAND3X1 U783 ( .IN1(n542), .IN2(n541), .IN3(n540), .OUT(n1158) );
  AOI22 U784 ( .IN1(n185), .IN2(n623), .IN3(Datain2[11]), .IN4(n746), .OUT(
        n545) );
  NAND3X1 U785 ( .IN1(n545), .IN2(n544), .IN3(n543), .OUT(n1160) );
  AOI22 U786 ( .IN1(n182), .IN2(n623), .IN3(Datain2[12]), .IN4(n746), .OUT(
        n548) );
  NAND3X1 U787 ( .IN1(n548), .IN2(n547), .IN3(n546), .OUT(n1161) );
  AOI22 U788 ( .IN1(n180), .IN2(n623), .IN3(Datain2[13]), .IN4(n746), .OUT(
        n551) );
  NAND3X1 U789 ( .IN1(n551), .IN2(n550), .IN3(n549), .OUT(n1162) );
  AOI22 U790 ( .IN1(n181), .IN2(n623), .IN3(Datain2[7]), .IN4(n746), .OUT(n554) );
  NAND3X1 U791 ( .IN1(n554), .IN2(n553), .IN3(n552), .OUT(n1156) );
  AOI22 U792 ( .IN1(Final_Exponent_reg[7]), .IN2(n623), .IN3(Datain2[14]), 
        .IN4(n746), .OUT(n557) );
  NAND3X1 U793 ( .IN1(n557), .IN2(n556), .IN3(n555), .OUT(n1164) );
  NOR2X1 U794 ( .IN1(Final_Exponent_reg[4]), .IN2(n180), .OUT(n559) );
  NOR2X1 U795 ( .IN1(n182), .IN2(Final_Exponent_reg[7]), .OUT(n558) );
  AOI22 U796 ( .IN1(n638), .IN2(n1115), .IN3(n733), .IN4(n710), .OUT(n570) );
  NOR2X1 U797 ( .IN1(Final_Exponent_reg[1]), .IN2(n184), .OUT(n563) );
  OAI21 U798 ( .IN1(n1112), .IN2(n628), .IN3(n568), .OUT(n569) );
  OAI21 U799 ( .IN1(n639), .IN2(n570), .IN3(n618), .OUT(n571) );
  AOI22 U800 ( .IN1(n653), .IN2(n1115), .IN3(n733), .IN4(n634), .OUT(n581) );
  NAND3X1 U801 ( .IN1(n220), .IN2(n196), .IN3(n639), .OUT(n576) );
  OAI21 U802 ( .IN1(n1112), .IN2(n708), .IN3(n579), .OUT(n580) );
  OAI21 U803 ( .IN1(n654), .IN2(n581), .IN3(n615), .OUT(n592) );
  NOR2X1 U804 ( .IN1(n650), .IN2(n648), .OUT(n585) );
  NOR2X1 U805 ( .IN1(n1112), .IN2(n650), .OUT(n584) );
  AOI22 U806 ( .IN1(n585), .IN2(n1115), .IN3(n584), .IN4(n583), .OUT(n591) );
  OAI21 U807 ( .IN1(n1112), .IN2(n636), .IN3(n588), .OUT(n589) );
  NOR2X1 U808 ( .IN1(n592), .IN2(n604), .OUT(n593) );
  NOR2X1 U809 ( .IN1(n657), .IN2(n660), .OUT(n597) );
  NOR2X1 U810 ( .IN1(n1112), .IN2(n660), .OUT(n596) );
  AOI22 U811 ( .IN1(n597), .IN2(n1115), .IN3(n596), .IN4(n595), .OUT(n612) );
  NOR2X1 U812 ( .IN1(n655), .IN2(n631), .OUT(n600) );
  NOR2X1 U813 ( .IN1(n1112), .IN2(n631), .OUT(n599) );
  AOI22 U814 ( .IN1(n600), .IN2(n1115), .IN3(n599), .IN4(n723), .OUT(n602) );
  NOR2X1 U815 ( .IN1(n604), .IN2(n603), .OUT(n605) );
  OAI21 U816 ( .IN1(n1097), .IN2(n607), .IN3(n667), .OUT(n608) );
  AOI21 U817 ( .IN1(n610), .IN2(n609), .IN3(n608), .OUT(n614) );
  NAND3X1 U818 ( .IN1(n733), .IN2(n629), .IN3(n630), .OUT(n613) );
  NAND3X1 U819 ( .IN1(n614), .IN2(n613), .IN3(n612), .OUT(n617) );
  NOR2X1 U820 ( .IN1(n617), .IN2(n616), .OUT(n620) );
  NAND3X1 U821 ( .IN1(n619), .IN2(n620), .IN3(n618), .OUT(C1_Z_0) );
  NAND3X1 U822 ( .IN1(n701), .IN2(n1191), .IN3(n1112), .OUT(n621) );
  NOR2X1 U823 ( .IN1(n712), .IN2(n621), .OUT(n622) );
  INVX4 U824 ( .IN(n622), .OUT(C2_Z_0) );
  AOI22 U825 ( .IN1(n183), .IN2(n623), .IN3(Datain2[10]), .IN4(n746), .OUT(
        n627) );
  NAND3X1 U826 ( .IN1(n627), .IN2(n626), .IN3(n625), .OUT(n1159) );
  AOI21 U827 ( .IN1(n637), .IN2(n674), .IN3(n1112), .OUT(n664) );
  AOI22 U828 ( .IN1(n641), .IN2(n640), .IN3(n639), .IN4(n638), .OUT(n642) );
  OAI21 U829 ( .IN1(n644), .IN2(n643), .IN3(n642), .OUT(n669) );
  NOR2X1 U830 ( .IN1(n755), .IN2(n669), .OUT(n645) );
  OAI21 U831 ( .IN1(n647), .IN2(n646), .IN3(n645), .OUT(n662) );
  AOI21 U832 ( .IN1(n662), .IN2(n1191), .IN3(n661), .OUT(n663) );
  AOI21 U833 ( .IN1(n677), .IN2(n664), .IN3(n663), .OUT(n796) );
  OAI21 U834 ( .IN1(n670), .IN2(n669), .IN3(n1115), .OUT(n671) );
  AOI21 U835 ( .IN1(n675), .IN2(n674), .IN3(n673), .OUT(n676) );
  OAI21 U836 ( .IN1(n677), .IN2(n1112), .IN3(n676), .OUT(n853) );
  AOI22 U837 ( .IN1(n1081), .IN2(n678), .IN3(n757), .IN4(n803), .OUT(n805) );
  OAI21 U838 ( .IN1(n265), .IN2(n1100), .IN3(n680), .OUT(n1117) );
  AOI22 U839 ( .IN1(Final_Mantissa_reg[10]), .IN2(n682), .IN3(n1115), .IN4(
        n681), .OUT(n683) );
  OAI21 U840 ( .IN1(n1112), .IN2(n727), .IN3(n683), .OUT(n684) );
  AOI22 U841 ( .IN1(Debug_reg[0]), .IN2(n1117), .IN3(n250), .IN4(n684), .OUT(
        n685) );
  AOI22 U842 ( .IN1(n751), .IN2(n688), .IN3(n687), .IN4(n686), .OUT(n1083) );
  AOI22 U843 ( .IN1(n692), .IN2(n691), .IN3(n690), .IN4(n689), .OUT(n1082) );
  AOI21 U844 ( .IN1(n750), .IN2(n194), .IN3(n693), .OUT(n694) );
  NOR2X1 U845 ( .IN1(n695), .IN2(n694), .OUT(n1087) );
  NOR2X1 U846 ( .IN1(n698), .IN2(n1097), .OUT(n703) );
  OAI21 U847 ( .IN1(n701), .IN2(n700), .IN3(n699), .OUT(n702) );
  AOI21 U848 ( .IN1(n1086), .IN2(n703), .IN3(n702), .OUT(n704) );
  OAI21 U849 ( .IN1(n706), .IN2(n705), .IN3(n704), .OUT(n1109) );
  NOR2X1 U850 ( .IN1(n1112), .IN2(n724), .OUT(n709) );
  NAND3X1 U851 ( .IN1(n709), .IN2(n708), .IN3(n726), .OUT(n711) );
  NOR2X1 U852 ( .IN1(n711), .IN2(n710), .OUT(n718) );
  NAND3X1 U853 ( .IN1(n714), .IN2(n713), .IN3(n712), .OUT(n715) );
  OAI21 U854 ( .IN1(n715), .IN2(n731), .IN3(n249), .OUT(n716) );
  AOI21 U855 ( .IN1(n718), .IN2(n717), .IN3(n716), .OUT(n719) );
  AOI22 U856 ( .IN1(n1115), .IN2(n722), .IN3(n721), .IN4(n720), .OUT(n1111) );
  AOI22 U857 ( .IN1(n253), .IN2(n224), .IN3(n258), .IN4(n825), .OUT(n734) );
  AOI22 U858 ( .IN1(n253), .IN2(n232), .IN3(n259), .IN4(n825), .OUT(n735) );
  AOI22 U859 ( .IN1(n253), .IN2(n227), .IN3(Final_Mantissa_reg[5]), .IN4(n825), 
        .OUT(n736) );
  AOI22 U860 ( .IN1(n253), .IN2(n225), .IN3(n260), .IN4(n825), .OUT(n737) );
  AOI22 U861 ( .IN1(n253), .IN2(n226), .IN3(n261), .IN4(n825), .OUT(n738) );
  AOI22 U862 ( .IN1(n253), .IN2(n228), .IN3(Final_Mantissa_reg[8]), .IN4(n825), 
        .OUT(n739) );
  AOI22 U863 ( .IN1(n253), .IN2(n231), .IN3(Final_Mantissa_reg[9]), .IN4(n825), 
        .OUT(n740) );
  AOI22 U864 ( .IN1(n253), .IN2(n185), .IN3(n182), .IN4(n825), .OUT(n741) );
  AOI22 U865 ( .IN1(n182), .IN2(n253), .IN3(n180), .IN4(n825), .OUT(
        ExcCheck_Datain_13__BAR) );
  AOI22 U866 ( .IN1(n180), .IN2(n253), .IN3(Final_Exponent_reg[7]), .IN4(n825), 
        .OUT(n742) );
  NOR2X1 U867 ( .IN1(n201), .IN2(Dataout_valid_BAR), .OUT(Dataout[0]) );
  NOR2X1 U868 ( .IN1(n203), .IN2(Dataout_valid_BAR), .OUT(Dataout[1]) );
  NOR2X1 U869 ( .IN1(n193), .IN2(Dataout_valid_BAR), .OUT(Dataout[2]) );
  NOR2X1 U870 ( .IN1(n222), .IN2(Dataout_valid_BAR), .OUT(Dataout[3]) );
  NOR2X1 U871 ( .IN1(n204), .IN2(Dataout_valid_BAR), .OUT(Dataout[4]) );
  NOR2X1 U872 ( .IN1(n195), .IN2(Dataout_valid_BAR), .OUT(Dataout[5]) );
  NOR2X1 U873 ( .IN1(n219), .IN2(Dataout_valid_BAR), .OUT(Dataout[6]) );
  NOR2X1 U874 ( .IN1(n233), .IN2(Dataout_valid_BAR), .OUT(Dataout[12]) );
  NOR2X1 U875 ( .IN1(n234), .IN2(Dataout_valid_BAR), .OUT(Dataout[13]) );
  NOR2X1 U876 ( .IN1(n235), .IN2(Dataout_valid_BAR), .OUT(Dataout[14]) );
  NOR2X1 U877 ( .IN1(Datain1[7]), .IN2(n936), .OUT(n760) );
  INVX1 U878 ( .IN(n775), .OUT(n758) );
  NOR2X1 U879 ( .IN1(Datain1[8]), .IN2(n935), .OUT(n773) );
  NOR2X1 U880 ( .IN1(n758), .IN2(n773), .OUT(n768) );
  INVX1 U881 ( .IN(n768), .OUT(n759) );
  AOI22 U882 ( .IN1(n760), .IN2(n768), .IN3(n759), .IN4(n767), .OUT(N152) );
  OAI21 U883 ( .IN1(n768), .IN2(n774), .IN3(n902), .OUT(N148) );
  OAI21 U884 ( .IN1(n760), .IN2(n773), .IN3(n775), .OUT(n762) );
  INVX1 U885 ( .IN(n762), .OUT(n761) );
  AOI22 U886 ( .IN1(Datain1[9]), .IN2(n763), .IN3(Datain2[9]), .IN4(n870), 
        .OUT(n777) );
  MUX2X1 U887 ( .IN1(n762), .IN2(n761), .S(n776), .OUT(n929) );
  NAND2X1 U888 ( .IN1(Datain2[9]), .IN2(n870), .OUT(n778) );
  AOI22 U889 ( .IN1(Datain1[9]), .IN2(n763), .IN3(n778), .IN4(n762), .OUT(n839) );
  INVX1 U890 ( .IN(n839), .OUT(n766) );
  INVX1 U891 ( .IN(Datain2[10]), .OUT(n764) );
  NOR2X1 U892 ( .IN1(Datain1[10]), .IN2(n764), .OUT(n878) );
  NAND2X1 U893 ( .IN1(Datain1[10]), .IN2(n764), .OUT(n880) );
  INVX1 U894 ( .IN(n880), .OUT(n765) );
  NOR2X1 U895 ( .IN1(n878), .IN2(n765), .OUT(n782) );
  MUX2X1 U896 ( .IN1(n766), .IN2(n839), .S(n782), .OUT(n913) );
  INVX1 U897 ( .IN(n913), .OUT(n772) );
  NAND2X1 U898 ( .IN1(n768), .IN2(n767), .OUT(n769) );
  NOR2X1 U899 ( .IN1(n264), .IN2(n769), .OUT(n1049) );
  AOI22 U900 ( .IN1(n929), .IN2(n770), .IN3(n1049), .IN4(n992), .OUT(N149) );
  NOR2X1 U901 ( .IN1(n992), .IN2(n770), .OUT(n771) );
  MUX2X1 U902 ( .IN1(n913), .IN2(n772), .S(n771), .OUT(N150) );
  NOR2X1 U903 ( .IN1(n179), .IN2(n252), .OUT(n1066) );
  AOI21 U904 ( .IN1(n775), .IN2(n774), .IN3(n773), .OUT(n779) );
  MUX2X1 U905 ( .IN1(n777), .IN2(n776), .S(n779), .OUT(n997) );
  NOR2X1 U906 ( .IN1(Datain2[9]), .IN2(n870), .OUT(n780) );
  OAI21 U907 ( .IN1(n780), .IN2(n779), .IN3(n778), .OUT(n879) );
  MUX2X1 U908 ( .IN1(n782), .IN2(n781), .S(n879), .OUT(n893) );
  NOR2X1 U909 ( .IN1(n264), .IN2(n902), .OUT(n982) );
  OAI21 U910 ( .IN1(n997), .IN2(n982), .IN3(n783), .OUT(N161) );
  MUX2X1 U911 ( .IN1(n784), .IN2(n893), .S(n783), .OUT(N162) );
  NAND2X1 U912 ( .IN1(StateMC[0]), .IN2(n198), .OUT(n785) );
  NOR2X1 U913 ( .IN1(StateMC[1]), .IN2(n785), .OUT(n826) );
  NAND3X1 U914 ( .IN1(StateMC[1]), .IN2(StateMC[2]), .IN3(n223), .OUT(n804) );
  OAI21 U915 ( .IN1(n253), .IN2(n825), .IN3(RSTn), .OUT(n1057) );
  NOR2X1 U916 ( .IN1(Exc_Ack), .IN2(n1057), .OUT(N274) );
  NAND2X1 U917 ( .IN1(StateMC[0]), .IN2(StateMC[2]), .OUT(n1056) );
  NOR2X1 U918 ( .IN1(StateMC[1]), .IN2(n1056), .OUT(n1081) );
  NOR2X1 U919 ( .IN1(n223), .IN2(n1100), .OUT(n1054) );
  INVX1 U920 ( .IN(Exc_value[0]), .OUT(n788) );
  INVX1 U921 ( .IN(Exc_value[2]), .OUT(n786) );
  AOI22 U922 ( .IN1(Exc_value[2]), .IN2(n788), .IN3(Exc_value[1]), .IN4(n786), 
        .OUT(n787) );
  OAI21 U923 ( .IN1(Exc_value[1]), .IN2(n788), .IN3(n787), .OUT(n789) );
  AOI22 U924 ( .IN1(n790), .IN2(n789), .IN3(StateMC[2]), .IN4(n223), .OUT(n791) );
  OAI21 U925 ( .IN1(n1081), .IN2(n792), .IN3(RSTn), .OUT(n958) );
  AOI22 U926 ( .IN1(n218), .IN2(n217), .IN3(exc_reg_0_), .IN4(n236), .OUT(n793) );
  AOI21 U927 ( .IN1(n217), .IN2(exc_reg_0_), .IN3(n793), .OUT(n828) );
  OAI21 U928 ( .IN1(n828), .IN2(n1108), .IN3(n794), .OUT(n812) );
  OAI21 U929 ( .IN1(n223), .IN2(n807), .IN3(n832), .OUT(n1106) );
  NOR2X1 U930 ( .IN1(n198), .IN2(StateMC[1]), .OUT(n1078) );
  AOI21 U931 ( .IN1(n796), .IN2(n1116), .IN3(n218), .OUT(n795) );
  NOR2X1 U932 ( .IN1(n835), .IN2(n795), .OUT(n852) );
  NOR2X1 U933 ( .IN1(n753), .IN2(n744), .OUT(n797) );
  AOI21 U934 ( .IN1(n796), .IN2(n797), .IN3(n217), .OUT(n848) );
  NAND2X1 U935 ( .IN1(n797), .IN2(n1112), .OUT(n799) );
  AOI22 U936 ( .IN1(n755), .IN2(n1191), .IN3(n743), .IN4(n229), .OUT(n798) );
  AOI21 U937 ( .IN1(n799), .IN2(exc_reg_0_), .IN3(n798), .OUT(n800) );
  MUX2X1 U938 ( .IN1(n852), .IN2(n848), .S(n853), .OUT(n802) );
  NAND2X1 U939 ( .IN1(n848), .IN2(n852), .OUT(n801) );
  NAND3X1 U940 ( .IN1(n1106), .IN2(n805), .IN3(n804), .OUT(n806) );
  OAI21 U941 ( .IN1(n812), .IN2(n806), .IN3(RSTn), .OUT(n965) );
  AOI22 U942 ( .IN1(StateMC[0]), .IN2(n809), .IN3(Exc_Ack), .IN4(n825), .OUT(
        n810) );
  NOR2X1 U943 ( .IN1(StateMC[2]), .IN2(n838), .OUT(n836) );
  NAND3X1 U944 ( .IN1(n810), .IN2(n1076), .IN3(n842), .OUT(n811) );
  OAI21 U945 ( .IN1(n812), .IN2(n811), .IN3(RSTn), .OUT(n1046) );
  NOR2X1 U946 ( .IN1(n223), .IN2(n199), .OUT(n845) );
  NOR2X1 U947 ( .IN1(n202), .IN2(Dataout_valid_BAR), .OUT(Dataout[10]) );
  NOR2X1 U948 ( .IN1(n230), .IN2(Dataout_valid_BAR), .OUT(Dataout[11]) );
  NOR2X1 U949 ( .IN1(n274), .IN2(Dataout_valid_BAR), .OUT(Dataout[15]) );
  NOR2X1 U950 ( .IN1(n220), .IN2(Dataout_valid_BAR), .OUT(Dataout[7]) );
  NOR2X1 U951 ( .IN1(n196), .IN2(Dataout_valid_BAR), .OUT(Dataout[8]) );
  NOR2X1 U952 ( .IN1(n205), .IN2(Dataout_valid_BAR), .OUT(Dataout[9]) );
  NAND2X1 U953 ( .IN1(Mode[0]), .IN2(n814), .OUT(n813) );
  NOR2X1 U954 ( .IN1(Mode[2]), .IN2(n813), .OUT(n819) );
  NOR2X1 U955 ( .IN1(Mode[2]), .IN2(n814), .OUT(n1192) );
  AOI22 U956 ( .IN1(StateMC[0]), .IN2(n819), .IN3(n1192), .IN4(Debug_reg[0]), 
        .OUT(n815) );
  AOI22 U957 ( .IN1(StateMC[1]), .IN2(n819), .IN3(n1192), .IN4(Debug_reg[1]), 
        .OUT(n816) );
  AOI22 U958 ( .IN1(StateMC[2]), .IN2(n819), .IN3(n1192), .IN4(Debug_reg[2]), 
        .OUT(n817) );
  NAND2X1 U959 ( .IN1(n1192), .IN2(Debug_reg[3]), .OUT(n818) );
  AOI21 U960 ( .IN1(Debug_valid_reg), .IN2(n1192), .IN3(n819), .OUT(n820) );
  AOI22 U961 ( .IN1(n253), .IN2(n184), .IN3(n183), .IN4(n825), .OUT(
        ExcCheck_Datain_10__BAR) );
  AOI22 U962 ( .IN1(n253), .IN2(n183), .IN3(n185), .IN4(n825), .OUT(n822) );
  AOI22 U963 ( .IN1(n253), .IN2(Op2_Mantissa_reg_7_), .IN3(n181), .IN4(n825), 
        .OUT(ExcCheck_Datain_7__BAR) );
  AOI22 U964 ( .IN1(n253), .IN2(n181), .IN3(n186), .IN4(n825), .OUT(n824) );
  AOI22 U965 ( .IN1(n253), .IN2(n186), .IN3(n184), .IN4(n825), .OUT(n827) );
  NOR2X1 U966 ( .IN1(Dataout_valid_BAR), .IN2(n828), .OUT(n829) );
  NOR2X1 U967 ( .IN1(n229), .IN2(n830), .OUT(Exc[0]) );
  NOR2X1 U968 ( .IN1(n218), .IN2(n830), .OUT(Exc[1]) );
  NOR2X1 U969 ( .IN1(n217), .IN2(n830), .OUT(Exc[2]) );
  NOR2X1 U970 ( .IN1(n265), .IN2(n831), .OUT(n1187) );
  NOR2X1 U971 ( .IN1(n214), .IN2(n1091), .OUT(N256) );
  NOR2X1 U972 ( .IN1(n213), .IN2(n1091), .OUT(N257) );
  NOR2X1 U973 ( .IN1(n212), .IN2(n1091), .OUT(N258) );
  NOR2X1 U974 ( .IN1(n211), .IN2(n1091), .OUT(N259) );
  NOR2X1 U975 ( .IN1(n210), .IN2(n1091), .OUT(N260) );
  NOR2X1 U976 ( .IN1(n209), .IN2(n1091), .OUT(N261) );
  NOR2X1 U977 ( .IN1(n208), .IN2(n1091), .OUT(N262) );
  NOR2X1 U978 ( .IN1(n207), .IN2(n1091), .OUT(N263) );
  NOR2X1 U979 ( .IN1(n265), .IN2(n1108), .OUT(n1094) );
  NAND3X1 U980 ( .IN1(RSTn), .IN2(n832), .IN3(n223), .OUT(n1090) );
  NAND3X1 U981 ( .IN1(n1090), .IN2(n1077), .IN3(n1091), .OUT(n833) );
  AOI22 U982 ( .IN1(Adder_dataout[8]), .IN2(n1094), .IN3(n206), .IN4(n833), 
        .OUT(n834) );
  OAI21 U983 ( .IN1(Data_valid), .IN2(n837), .IN3(n1090), .OUT(n859) );
  OAI21 U984 ( .IN1(n878), .IN2(n839), .IN3(n880), .OUT(n916) );
  NAND2X1 U985 ( .IN1(Datain2[11]), .IN2(n892), .OUT(n881) );
  AOI22 U986 ( .IN1(Datain1[11]), .IN2(n933), .IN3(n916), .IN4(n881), .OUT(
        n928) );
  NAND2X1 U987 ( .IN1(Datain1[12]), .IN2(n932), .OUT(n883) );
  INVX1 U988 ( .IN(Datain1[12]), .OUT(n884) );
  AOI22 U989 ( .IN1(n928), .IN2(n883), .IN3(Datain2[12]), .IN4(n884), .OUT(
        n924) );
  INVX1 U990 ( .IN(Datain1[13]), .OUT(n911) );
  NAND2X1 U991 ( .IN1(Datain2[13]), .IN2(n911), .OUT(n910) );
  AOI22 U992 ( .IN1(n924), .IN2(n910), .IN3(Datain1[13]), .IN4(n840), .OUT(
        n920) );
  AOI22 U993 ( .IN1(n920), .IN2(n841), .IN3(Datain2[14]), .IN4(n885), .OUT(
        n844) );
  NOR2X1 U994 ( .IN1(n265), .IN2(n842), .OUT(n843) );
  AOI21 U995 ( .IN1(RSTn), .IN2(n845), .IN3(N274), .OUT(n846) );
  NAND3X1 U996 ( .IN1(n846), .IN2(n1090), .IN3(n1096), .OUT(n850) );
  INVX1 U997 ( .IN(Exc_Ack), .OUT(n847) );
  NOR2X1 U998 ( .IN1(n847), .IN2(n1057), .OUT(n854) );
  AOI22 U999 ( .IN1(n848), .IN2(n250), .IN3(n854), .IN4(Exc_value[2]), .OUT(
        n849) );
  OAI21 U1000 ( .IN1(n217), .IN2(n856), .IN3(n849), .OUT(n1163) );
  AOI22 U1001 ( .IN1(Exc_value[1]), .IN2(n854), .IN3(n236), .IN4(n850), .OUT(
        n851) );
  OAI21 U1002 ( .IN1(n852), .IN2(n1193), .IN3(n851), .OUT(n1155) );
  AOI22 U1003 ( .IN1(Exc_value[0]), .IN2(n854), .IN3(n250), .IN4(n853), .OUT(
        n855) );
  OAI21 U1004 ( .IN1(n856), .IN2(n229), .IN3(n855), .OUT(n1154) );
  AOI21 U1005 ( .IN1(n857), .IN2(Adder_valid), .IN3(n254), .OUT(n858) );
  AOI21 U1006 ( .IN1(RSTn), .IN2(n860), .IN3(n859), .OUT(n877) );
  AOI22 U1007 ( .IN1(n745), .IN2(Datain2[15]), .IN3(n746), .IN4(Datain1[15]), 
        .OUT(n861) );
  OAI21 U1008 ( .IN1(n215), .IN2(n255), .IN3(n861), .OUT(n1152) );
  AOI22 U1009 ( .IN1(n745), .IN2(Datain1[0]), .IN3(n746), .IN4(Datain2[0]), 
        .OUT(n862) );
  OAI21 U1010 ( .IN1(n255), .IN2(n214), .IN3(n862), .OUT(n1151) );
  AOI22 U1011 ( .IN1(n745), .IN2(Datain1[1]), .IN3(n746), .IN4(Datain2[1]), 
        .OUT(n863) );
  OAI21 U1012 ( .IN1(n255), .IN2(n213), .IN3(n863), .OUT(n1150) );
  AOI22 U1013 ( .IN1(n745), .IN2(Datain1[2]), .IN3(n746), .IN4(Datain2[2]), 
        .OUT(n864) );
  OAI21 U1014 ( .IN1(n255), .IN2(n212), .IN3(n864), .OUT(n1149) );
  AOI22 U1015 ( .IN1(n745), .IN2(Datain1[3]), .IN3(n746), .IN4(Datain2[3]), 
        .OUT(n865) );
  OAI21 U1016 ( .IN1(n255), .IN2(n211), .IN3(n865), .OUT(n1148) );
  AOI22 U1017 ( .IN1(n745), .IN2(Datain1[4]), .IN3(n746), .IN4(Datain2[4]), 
        .OUT(n866) );
  OAI21 U1018 ( .IN1(n255), .IN2(n210), .IN3(n866), .OUT(n1147) );
  AOI22 U1019 ( .IN1(n745), .IN2(n256), .IN3(n746), .IN4(Datain2[5]), .OUT(
        n867) );
  OAI21 U1020 ( .IN1(n255), .IN2(n209), .IN3(n867), .OUT(n1146) );
  AOI22 U1021 ( .IN1(n745), .IN2(n257), .IN3(n746), .IN4(Datain2[6]), .OUT(
        n868) );
  OAI21 U1022 ( .IN1(n255), .IN2(n208), .IN3(n868), .OUT(n1145) );
  NOR2X1 U1023 ( .IN1(Datain1[13]), .IN2(Datain1[10]), .OUT(n869) );
  NAND3X1 U1024 ( .IN1(n870), .IN2(n885), .IN3(n869), .OUT(n873) );
  NOR2X1 U1025 ( .IN1(Datain1[8]), .IN2(Datain1[7]), .OUT(n871) );
  NAND3X1 U1026 ( .IN1(n884), .IN2(n871), .IN3(n892), .OUT(n872) );
  NOR2X1 U1027 ( .IN1(n873), .IN2(n872), .OUT(n943) );
  OAI21 U1028 ( .IN1(n1071), .IN2(n943), .IN3(n1073), .OUT(n874) );
  OAI21 U1029 ( .IN1(n255), .IN2(n207), .IN3(n875), .OUT(n1144) );
  AOI22 U1030 ( .IN1(n745), .IN2(Datain1[15]), .IN3(n746), .IN4(Datain2[15]), 
        .OUT(n876) );
  OAI21 U1031 ( .IN1(n191), .IN2(n255), .IN3(n876), .OUT(n1143) );
  OAI21 U1032 ( .IN1(Datain1[12]), .IN2(n932), .IN3(n883), .OUT(n909) );
  NOR2X1 U1033 ( .IN1(Datain2[11]), .IN2(n892), .OUT(n882) );
  AOI21 U1034 ( .IN1(n880), .IN2(n879), .IN3(n878), .OUT(n895) );
  OAI21 U1035 ( .IN1(n882), .IN2(n895), .IN3(n881), .OUT(n900) );
  AOI22 U1036 ( .IN1(Datain2[12]), .IN2(n884), .IN3(n883), .IN4(n900), .OUT(
        n888) );
  AOI22 U1037 ( .IN1(Datain1[14]), .IN2(n886), .IN3(Datain2[14]), .IN4(n885), 
        .OUT(n919) );
  NOR2X1 U1038 ( .IN1(Datain2[13]), .IN2(n911), .OUT(n887) );
  MUX2X1 U1039 ( .IN1(n919), .IN2(n888), .S(n887), .OUT(n889) );
  MUX2X1 U1040 ( .IN1(n891), .IN2(n890), .S(n910), .OUT(n897) );
  AOI22 U1041 ( .IN1(Datain1[11]), .IN2(n933), .IN3(Datain2[11]), .IN4(n892), 
        .OUT(n912) );
  AOI21 U1042 ( .IN1(n912), .IN2(n895), .IN3(n893), .OUT(n894) );
  OAI21 U1043 ( .IN1(n912), .IN2(n895), .IN3(n894), .OUT(n896) );
  NOR2X1 U1044 ( .IN1(n897), .IN2(n896), .OUT(n898) );
  OAI21 U1045 ( .IN1(n909), .IN2(n900), .IN3(n898), .OUT(n899) );
  AOI21 U1046 ( .IN1(n909), .IN2(n900), .IN3(n899), .OUT(n946) );
  INVX1 U1047 ( .IN(n946), .OUT(n901) );
  NOR2X1 U1048 ( .IN1(n901), .IN2(n1014), .OUT(n987) );
  INVX1 U1049 ( .IN(Datain1[3]), .OUT(n996) );
  NOR2X1 U1050 ( .IN1(n179), .IN2(N156), .OUT(n1074) );
  INVX1 U1051 ( .IN(Datain1[1]), .OUT(n903) );
  AOI22 U1052 ( .IN1(n1066), .IN2(n996), .IN3(n1074), .IN4(n903), .OUT(n904)
         );
  OAI21 U1053 ( .IN1(Datain1[2]), .IN2(n980), .IN3(n904), .OUT(n907) );
  NAND2X1 U1054 ( .IN1(n982), .IN2(Datain1[4]), .OUT(n905) );
  OAI21 U1055 ( .IN1(n979), .IN2(n980), .IN3(n905), .OUT(n906) );
  AOI21 U1056 ( .IN1(n1074), .IN2(n256), .IN3(n906), .OUT(n1030) );
  AOI22 U1057 ( .IN1(n997), .IN2(n907), .IN3(n1030), .IN4(n984), .OUT(n908) );
  AOI22 U1058 ( .IN1(n987), .IN2(n908), .IN3(n224), .IN4(n1051), .OUT(n956) );
  OAI21 U1059 ( .IN1(Datain2[13]), .IN2(n911), .IN3(n910), .OUT(n923) );
  AOI21 U1060 ( .IN1(n916), .IN2(n915), .IN3(n913), .OUT(n914) );
  OAI21 U1061 ( .IN1(n916), .IN2(n915), .IN3(n914), .OUT(n917) );
  AOI21 U1062 ( .IN1(n920), .IN2(n919), .IN3(n917), .OUT(n918) );
  OAI21 U1063 ( .IN1(n920), .IN2(n919), .IN3(n918), .OUT(n921) );
  AOI21 U1064 ( .IN1(n924), .IN2(n923), .IN3(n921), .OUT(n922) );
  OAI21 U1065 ( .IN1(n924), .IN2(n923), .IN3(n922), .OUT(n925) );
  AOI21 U1066 ( .IN1(n928), .IN2(n927), .IN3(n925), .OUT(n926) );
  OAI21 U1067 ( .IN1(n928), .IN2(n927), .IN3(n926), .OUT(n994) );
  NOR2X1 U1068 ( .IN1(n929), .IN2(n994), .OUT(n1010) );
  INVX1 U1069 ( .IN(Datain2[6]), .OUT(n957) );
  INVX1 U1070 ( .IN(Datain2[4]), .OUT(n930) );
  AOI22 U1071 ( .IN1(N168), .IN2(n957), .IN3(n930), .IN4(n251), .OUT(n1020) );
  NOR2X1 U1072 ( .IN1(n179), .IN2(N168), .OUT(n962) );
  AOI22 U1073 ( .IN1(n179), .IN2(n1020), .IN3(Datain2[5]), .IN4(n962), .OUT(
        n942) );
  NOR2X1 U1074 ( .IN1(Datain2[14]), .IN2(Datain2[13]), .OUT(n931) );
  NAND3X1 U1075 ( .IN1(n933), .IN2(n932), .IN3(n931), .OUT(n938) );
  NOR2X1 U1076 ( .IN1(Datain2[10]), .IN2(Datain2[9]), .OUT(n934) );
  NAND3X1 U1077 ( .IN1(n936), .IN2(n935), .IN3(n934), .OUT(n937) );
  NOR2X1 U1078 ( .IN1(n938), .IN2(n937), .OUT(n1009) );
  NOR2X1 U1079 ( .IN1(n1009), .IN2(n1071), .OUT(n1052) );
  NOR2X1 U1080 ( .IN1(N168), .IN2(Datain2[5]), .OUT(n959) );
  AOI22 U1081 ( .IN1(N168), .IN2(Datain2[6]), .IN3(Datain2[4]), .IN4(n1049), 
        .OUT(n939) );
  OAI21 U1082 ( .IN1(n179), .IN2(n959), .IN3(n939), .OUT(n940) );
  OAI21 U1083 ( .IN1(n942), .IN2(n1002), .IN3(n941), .OUT(n1032) );
  NOR2X1 U1084 ( .IN1(n943), .IN2(n1073), .OUT(n947) );
  NAND2X1 U1085 ( .IN1(n946), .IN2(n947), .OUT(n995) );
  NOR2X1 U1086 ( .IN1(n997), .IN2(n995), .OUT(n990) );
  NOR2X1 U1087 ( .IN1(n264), .IN2(n257), .OUT(n945) );
  AOI22 U1088 ( .IN1(Datain1[4]), .IN2(n982), .IN3(n256), .IN4(N366), .OUT(
        n944) );
  OAI21 U1089 ( .IN1(n252), .IN2(n945), .IN3(n944), .OUT(n1029) );
  AOI22 U1090 ( .IN1(n1010), .IN2(n1032), .IN3(n990), .IN4(n1029), .OUT(n955)
         );
  INVX1 U1091 ( .IN(Datain1[2]), .OUT(n970) );
  NOR2X1 U1092 ( .IN1(n992), .IN2(n994), .OUT(n1067) );
  NOR2X1 U1093 ( .IN1(N168), .IN2(n1019), .OUT(n967) );
  NOR2X1 U1094 ( .IN1(n251), .IN2(n1019), .OUT(n1000) );
  AOI22 U1095 ( .IN1(n967), .IN2(Datain2[0]), .IN3(n1000), .IN4(Datain2[2]), 
        .OUT(n948) );
  OAI21 U1096 ( .IN1(n949), .IN2(n970), .IN3(n948), .OUT(n953) );
  AOI22 U1097 ( .IN1(Datain1[3]), .IN2(n1001), .IN3(Datain2[3]), .IN4(n1000), 
        .OUT(n952) );
  NOR2X1 U1098 ( .IN1(N156), .IN2(n950), .OUT(n1044) );
  AOI22 U1099 ( .IN1(n1044), .IN2(Datain1[1]), .IN3(n967), .IN4(Datain2[1]), 
        .OUT(n951) );
  AOI22 U1100 ( .IN1(n179), .IN2(n953), .IN3(n966), .IN4(N366), .OUT(n954) );
  NAND3X1 U1101 ( .IN1(n956), .IN2(n955), .IN3(n954), .OUT(n1142) );
  NAND2X1 U1102 ( .IN1(Datain2[5]), .IN2(n1049), .OUT(n964) );
  NOR2X1 U1103 ( .IN1(n1071), .IN2(n957), .OUT(n961) );
  NOR2X1 U1104 ( .IN1(n959), .IN2(N366), .OUT(n960) );
  AOI22 U1105 ( .IN1(n962), .IN2(n961), .IN3(n1052), .IN4(n960), .OUT(n963) );
  OAI21 U1106 ( .IN1(n1002), .IN2(n964), .IN3(n963), .OUT(n1035) );
  AOI22 U1107 ( .IN1(n179), .IN2(n966), .IN3(n1010), .IN4(n1035), .OUT(n978)
         );
  AOI22 U1108 ( .IN1(n1001), .IN2(Datain1[4]), .IN3(n1000), .IN4(Datain2[4]), 
        .OUT(n969) );
  AOI22 U1109 ( .IN1(n1044), .IN2(Datain1[2]), .IN3(n967), .IN4(Datain2[2]), 
        .OUT(n968) );
  INVX1 U1110 ( .IN(Datain1[4]), .OUT(n981) );
  AOI22 U1111 ( .IN1(n1066), .IN2(n981), .IN3(n1074), .IN4(n970), .OUT(n971)
         );
  OAI21 U1112 ( .IN1(Datain1[3]), .IN2(n980), .IN3(n971), .OUT(n972) );
  AOI22 U1113 ( .IN1(n1074), .IN2(n257), .IN3(n256), .IN4(n982), .OUT(n1036)
         );
  AOI22 U1114 ( .IN1(n997), .IN2(n972), .IN3(n1036), .IN4(n984), .OUT(n974) );
  AOI22 U1115 ( .IN1(n179), .IN2(n256), .IN3(n1074), .IN4(n257), .OUT(n973) );
  AOI22 U1116 ( .IN1(n987), .IN2(n974), .IN3(n990), .IN4(n1039), .OUT(n975) );
  OAI21 U1117 ( .IN1(n1028), .IN2(add_x_35_A_4_), .IN3(n975), .OUT(n976) );
  AOI21 U1118 ( .IN1(n264), .IN2(n1007), .IN3(n976), .OUT(n977) );
  NOR2X1 U1119 ( .IN1(N156), .IN2(n979), .OUT(n991) );
  AOI22 U1120 ( .IN1(n1066), .IN2(n1015), .IN3(n1016), .IN4(n981), .OUT(n986)
         );
  AOI22 U1121 ( .IN1(n1074), .IN2(n996), .IN3(n984), .IN4(n983), .OUT(n985) );
  NAND3X1 U1122 ( .IN1(n987), .IN2(n986), .IN3(n985), .OUT(n988) );
  OAI21 U1123 ( .IN1(n1028), .IN2(add_x_35_A_5_), .IN3(n988), .OUT(n989) );
  AOI21 U1124 ( .IN1(n991), .IN2(n990), .IN3(n989), .OUT(n1013) );
  OAI21 U1125 ( .IN1(n992), .IN2(Datain2[3]), .IN3(n1052), .OUT(n993) );
  NOR2X1 U1126 ( .IN1(n994), .IN2(n993), .OUT(n999) );
  AOI21 U1127 ( .IN1(n997), .IN2(n996), .IN3(n995), .OUT(n998) );
  AOI22 U1128 ( .IN1(n999), .IN2(n251), .IN3(n998), .IN4(n252), .OUT(n1006) );
  AOI22 U1129 ( .IN1(n1001), .IN2(n256), .IN3(n1000), .IN4(Datain2[5]), .OUT(
        n1005) );
  NAND3X1 U1130 ( .IN1(Datain2[3]), .IN2(n1003), .IN3(n1072), .OUT(n1004) );
  NAND3X1 U1131 ( .IN1(n1006), .IN2(n1005), .IN3(n1004), .OUT(n1017) );
  AOI22 U1132 ( .IN1(n179), .IN2(n1007), .IN3(n1017), .IN4(n264), .OUT(n1012)
         );
  NAND2X1 U1133 ( .IN1(n745), .IN2(Datain2[6]), .OUT(n1008) );
  AOI21 U1134 ( .IN1(n1009), .IN2(N366), .IN3(n1008), .OUT(n1043) );
  NAND3X1 U1135 ( .IN1(n1010), .IN2(n1043), .IN3(n251), .OUT(n1011) );
  NAND3X1 U1136 ( .IN1(n1013), .IN2(n1012), .IN3(n1011), .OUT(n1140) );
  NOR2X1 U1137 ( .IN1(n1065), .IN2(n1014), .OUT(n1038) );
  AOI22 U1138 ( .IN1(N156), .IN2(n257), .IN3(Datain1[4]), .IN4(n252), .OUT(
        n1018) );
  AOI22 U1139 ( .IN1(n1016), .IN2(n1015), .IN3(n1018), .IN4(n264), .OUT(n1026)
         );
  INVX1 U1140 ( .IN(n1017), .OUT(n1024) );
  INVX1 U1141 ( .IN(n1019), .OUT(n1021) );
  AOI22 U1142 ( .IN1(n1040), .IN2(n1022), .IN3(n1021), .IN4(n1020), .OUT(n1023) );
  AOI22 U1143 ( .IN1(n179), .IN2(n1024), .IN3(n1023), .IN4(n264), .OUT(n1025)
         );
  AOI21 U1144 ( .IN1(n1038), .IN2(n1026), .IN3(n1025), .OUT(n1027) );
  OAI21 U1145 ( .IN1(n1028), .IN2(add_x_35_A_6_), .IN3(n1027), .OUT(n1139) );
  AOI22 U1146 ( .IN1(n1040), .IN2(n1029), .IN3(n1051), .IN4(n226), .OUT(n1034)
         );
  AOI22 U1147 ( .IN1(n1067), .IN2(n1032), .IN3(n1038), .IN4(n1031), .OUT(n1033) );
  AOI22 U1148 ( .IN1(n1067), .IN2(n1035), .IN3(n1051), .IN4(n228), .OUT(n1042)
         );
  AOI22 U1149 ( .IN1(n1040), .IN2(n1039), .IN3(n1038), .IN4(n1037), .OUT(n1041) );
  AOI21 U1150 ( .IN1(n1052), .IN2(N366), .IN3(n1043), .OUT(n1048) );
  AOI21 U1151 ( .IN1(n1051), .IN2(n231), .IN3(n1044), .OUT(n1045) );
  OAI21 U1152 ( .IN1(n1048), .IN2(n1047), .IN3(n1045), .OUT(n1136) );
  NAND2X1 U1153 ( .IN1(n1067), .IN2(n1049), .OUT(n1050) );
  AOI22 U1154 ( .IN1(n1061), .IN2(n1052), .IN3(Op2_Mantissa_reg_7_), .IN4(
        n1051), .OUT(n1053) );
  NOR2X1 U1155 ( .IN1(n200), .IN2(n238), .OUT(n1118) );
  MUX2X1 U1156 ( .IN1(add_x_35_A_2_), .IN2(n237), .S(n1118), .OUT(n1060) );
  OAI21 U1157 ( .IN1(n756), .IN2(Adder_ack), .IN3(n1054), .OUT(n1055) );
  NAND3X1 U1158 ( .IN1(n1090), .IN2(n1193), .IN3(n1057), .OUT(n1058) );
  AOI21 U1159 ( .IN1(RSTn), .IN2(n1059), .IN3(n1058), .OUT(n1068) );
  AOI22 U1160 ( .IN1(n1060), .IN2(n1070), .IN3(n237), .IN4(n1069), .OUT(n1064)
         );
  NOR2X1 U1161 ( .IN1(n1061), .IN2(n1071), .OUT(n1062) );
  AOI22 U1162 ( .IN1(n746), .IN2(N434), .IN3(N380), .IN4(n1062), .OUT(n1063)
         );
  AOI21 U1163 ( .IN1(n1087), .IN2(n1086), .IN3(n1085), .OUT(n1089) );
  NOR2X1 U1164 ( .IN1(n1190), .IN2(n250), .OUT(n1093) );
  NAND3X1 U1165 ( .IN1(n1093), .IN2(n1092), .IN3(n1091), .OUT(n1095) );
  AOI21 U1166 ( .IN1(n215), .IN2(n1097), .IN3(n191), .OUT(n1098) );
  NOR2X1 U1167 ( .IN1(n753), .IN2(n1098), .OUT(n1103) );
  NOR2X1 U1168 ( .IN1(n277), .IN2(n1099), .OUT(n1101) );
  AOI22 U1169 ( .IN1(RSTn), .IN2(n1101), .IN3(n1117), .IN4(n241), .OUT(n1102)
         );
  OAI21 U1170 ( .IN1(n1193), .IN2(n1103), .IN3(n1102), .OUT(n1122) );
  AOI22 U1171 ( .IN1(n749), .IN2(n751), .IN3(n750), .IN4(n754), .OUT(n1105) );
  NAND3X1 U1172 ( .IN1(n1106), .IN2(n1105), .IN3(n1104), .OUT(n1107) );
  AOI22 U1173 ( .IN1(n250), .IN2(n1109), .IN3(Debug_reg[2]), .IN4(n1117), 
        .OUT(n1110) );
  OAI21 U1174 ( .IN1(n752), .IN2(n1112), .IN3(n1111), .OUT(n1113) );
  AOI22 U1175 ( .IN1(n250), .IN2(n1113), .IN3(Debug_reg[1]), .IN4(n1117), 
        .OUT(n1114) );
  NOR2X1 U1176 ( .IN1(n224), .IN2(n1185), .OUT(n1182) );
  NOR2X1 U1177 ( .IN1(n227), .IN2(n1179), .OUT(n1176) );
  NAND2X1 U1178 ( .IN1(add_x_35_A_6_), .IN2(n1176), .OUT(n1173) );
  NOR2X1 U1179 ( .IN1(n226), .IN2(n1173), .OUT(n1170) );
  NOR2X1 U1180 ( .IN1(n231), .IN2(n1167), .OUT(n1120) );
  AOI21 U1181 ( .IN1(n1120), .IN2(n239), .IN3(n1119), .OUT(n114) );
  NOR2X1 U1182 ( .IN1(n1120), .IN2(n756), .OUT(n1166) );
  OAI21 U1183 ( .IN1(Op2_Mantissa_reg_7_), .IN2(n1166), .IN3(n254), .OUT(n1121) );
  AOI21 U1184 ( .IN1(Op2_Mantissa_reg_7_), .IN2(n1166), .IN3(n1121), .OUT(n113) );
  OAI21 U1185 ( .IN1(add_x_35_A_9_), .IN2(n1169), .IN3(n254), .OUT(n1168) );
  AOI21 U1186 ( .IN1(add_x_35_A_9_), .IN2(n1169), .IN3(n1168), .OUT(n112) );
  NOR2X1 U1187 ( .IN1(n1170), .IN2(n756), .OUT(n1172) );
  OAI21 U1188 ( .IN1(n1172), .IN2(n228), .IN3(n254), .OUT(n1171) );
  AOI21 U1189 ( .IN1(n1172), .IN2(n228), .IN3(n1171), .OUT(n111) );
  OAI21 U1190 ( .IN1(add_x_35_A_7_), .IN2(n1175), .IN3(n254), .OUT(n1174) );
  AOI21 U1191 ( .IN1(add_x_35_A_7_), .IN2(n1175), .IN3(n1174), .OUT(n110) );
  NOR2X1 U1192 ( .IN1(n1176), .IN2(n756), .OUT(n1178) );
  OAI21 U1193 ( .IN1(n1178), .IN2(n225), .IN3(n254), .OUT(n1177) );
  AOI21 U1194 ( .IN1(n1178), .IN2(n225), .IN3(n1177), .OUT(n109) );
  OAI21 U1195 ( .IN1(add_x_35_A_5_), .IN2(n1181), .IN3(n254), .OUT(n1180) );
  AOI21 U1196 ( .IN1(add_x_35_A_5_), .IN2(n1181), .IN3(n1180), .OUT(n108) );
  NOR2X1 U1197 ( .IN1(n1182), .IN2(n756), .OUT(n1184) );
  OAI21 U1198 ( .IN1(n1184), .IN2(n232), .IN3(n254), .OUT(n1183) );
  AOI21 U1199 ( .IN1(n1184), .IN2(n232), .IN3(n1183), .OUT(n107) );
  OAI21 U1200 ( .IN1(add_x_35_A_3_), .IN2(n1189), .IN3(n254), .OUT(n1188) );
  AOI21 U1201 ( .IN1(add_x_35_A_3_), .IN2(n1189), .IN3(n1188), .OUT(n106) );
  MUX2X1 U1202 ( .IN1(n1200), .IN2(n1201), .S(n252), .OUT(n1194) );
  MUX2X1 U1203 ( .IN1(n1202), .IN2(n1203), .S(n252), .OUT(n1195) );
  MUX2X1 U1204 ( .IN1(n1204), .IN2(n1205), .S(n252), .OUT(n1196) );
  MUX2X1 U1205 ( .IN1(n1206), .IN2(n1207), .S(n252), .OUT(n1197) );
  MUX2X1 U1206 ( .IN1(n1194), .IN2(n1195), .S(N149), .OUT(n1198) );
  MUX2X1 U1207 ( .IN1(n1196), .IN2(n1197), .S(N149), .OUT(n1199) );
  MUX2X1 U1208 ( .IN1(n1198), .IN2(n1199), .S(N150), .OUT(N380) );
  MUX2X1 U1209 ( .IN1(Datain2[0]), .IN2(Datain2[1]), .S(n179), .OUT(n1200) );
  MUX2X1 U1210 ( .IN1(Datain2[2]), .IN2(Datain2[3]), .S(n179), .OUT(n1201) );
  MUX2X1 U1211 ( .IN1(Datain2[4]), .IN2(Datain2[5]), .S(n179), .OUT(n1202) );
  MUX2X1 U1212 ( .IN1(Datain2[6]), .IN2(Datain2[7]), .S(n179), .OUT(n1203) );
  MUX2X1 U1213 ( .IN1(Datain2[8]), .IN2(Datain2[9]), .S(n179), .OUT(n1204) );
  MUX2X1 U1214 ( .IN1(Datain2[10]), .IN2(Datain2[11]), .S(n179), .OUT(n1205)
         );
  MUX2X1 U1215 ( .IN1(Datain2[12]), .IN2(Datain2[13]), .S(n179), .OUT(n1206)
         );
  MUX2X1 U1216 ( .IN1(Datain2[14]), .IN2(Datain2[15]), .S(n179), .OUT(n1207)
         );
  MUX2X1 U1217 ( .IN1(n1218), .IN2(n1219), .S(n251), .OUT(n1208) );
  MUX2X1 U1218 ( .IN1(n1220), .IN2(n1221), .S(n251), .OUT(n1209) );
  MUX2X1 U1219 ( .IN1(n1222), .IN2(n1223), .S(n251), .OUT(n1210) );
  MUX2X1 U1220 ( .IN1(n1224), .IN2(n1225), .S(n251), .OUT(n1211) );
  MUX2X1 U1221 ( .IN1(n1208), .IN2(n1209), .S(N161), .OUT(n1212) );
  MUX2X1 U1222 ( .IN1(n1210), .IN2(n1211), .S(N161), .OUT(n1213) );
  MUX2X1 U1223 ( .IN1(n1212), .IN2(n1213), .S(N162), .OUT(N434) );
  MUX2X1 U1224 ( .IN1(Datain1[0]), .IN2(Datain1[1]), .S(N366), .OUT(n1214) );
  MUX2X1 U1225 ( .IN1(Datain1[2]), .IN2(Datain1[3]), .S(N366), .OUT(n1215) );
  MUX2X1 U1226 ( .IN1(Datain1[4]), .IN2(n256), .S(n264), .OUT(n1216) );
  MUX2X1 U1227 ( .IN1(n257), .IN2(Datain1[7]), .S(N366), .OUT(n1217) );
  MUX2X1 U1228 ( .IN1(Datain1[0]), .IN2(Datain1[1]), .S(n179), .OUT(n1218) );
  MUX2X1 U1229 ( .IN1(Datain1[2]), .IN2(Datain1[3]), .S(n179), .OUT(n1219) );
  MUX2X1 U1230 ( .IN1(Datain1[4]), .IN2(n256), .S(n179), .OUT(n1220) );
  MUX2X1 U1231 ( .IN1(n257), .IN2(Datain1[7]), .S(n179), .OUT(n1221) );
  MUX2X1 U1232 ( .IN1(Datain1[8]), .IN2(Datain1[9]), .S(n179), .OUT(n1222) );
  MUX2X1 U1233 ( .IN1(Datain1[10]), .IN2(Datain1[11]), .S(n179), .OUT(n1223)
         );
  MUX2X1 U1234 ( .IN1(Datain1[12]), .IN2(Datain1[13]), .S(n179), .OUT(n1224)
         );
  MUX2X1 U1235 ( .IN1(Datain1[14]), .IN2(Datain1[15]), .S(n179), .OUT(n1225)
         );
endmodule


module Mul_cntrl ( CLK, RSTn, Datain1, Datain2, Data_valid, Dataout, 
        Dataout_valid, Exc, Mode, Debug, Multi_datain1, Multi_datain2, 
        Multi_dataout, Multi_ack, ExcCheck_valid, ExcCheck_Datain, Exc_value, 
        Multi_valid_BAR, Exc_Ack_BAR );
  input [15:0] Datain1;
  input [15:0] Datain2;
  output [15:0] Dataout;
  output [2:0] Exc;
  input [2:0] Mode;
  output [4:0] Debug;
  output [7:0] Multi_datain1;
  output [7:0] Multi_datain2;
  input [15:0] Multi_dataout;
  output [15:0] ExcCheck_Datain;
  input [2:0] Exc_value;
  input CLK, RSTn, Data_valid, Multi_ack, Exc_Ack_BAR;
  output Dataout_valid, ExcCheck_valid, Multi_valid_BAR;
  wire   Debug_valid_reg, Final_Sign_reg, G_reg, T_reg, N89, N90, N384, N385,
         N386, N387, N388, N389, N390, N391, N392, C276_DATA3_0, C276_DATA3_1,
         C276_DATA3_2, C276_DATA3_3, C276_DATA3_8, n64, n94, n96, n124, n125,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n144, n145, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n213, n214, n215, n667, n703, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, C1_Z_3, C1_Z_1, C1_Z_0,
         RSOP_428_C1_Z_0, DP_OP_357J3_124_4634_n29, DP_OP_357J3_124_4634_n28,
         DP_OP_357J3_124_4634_n27, DP_OP_357J3_124_4634_n26,
         DP_OP_357J3_124_4634_n25, DP_OP_357J3_124_4634_n24,
         DP_OP_357J3_124_4634_n23, DP_OP_357J3_124_4634_n22,
         DP_OP_357J3_124_4634_n21, DP_OP_357J3_124_4634_n20,
         DP_OP_357J3_124_4634_n19, DP_OP_357J3_124_4634_n18,
         DP_OP_357J3_124_4634_n17, DP_OP_357J3_124_4634_n15,
         DP_OP_357J3_124_4634_n13, DP_OP_357J3_124_4634_n12,
         DP_OP_357J3_124_4634_n11, DP_OP_357J3_124_4634_n10,
         DP_OP_357J3_124_4634_n9, DP_OP_357J3_124_4634_n8,
         DP_OP_357J3_124_4634_n7, DP_OP_357J3_124_4634_n6,
         DP_OP_357J3_124_4634_n5, DP_OP_357J3_124_4634_n4,
         DP_OP_357J3_124_4634_n3, DP_OP_357J3_124_4634_n2,
         DP_OP_357J3_124_4634_n1, DP_OP_433J3_126_901_n30,
         DP_OP_433J3_126_901_n29, DP_OP_433J3_126_901_n28,
         DP_OP_433J3_126_901_n23, DP_OP_433J3_126_901_n21,
         DP_OP_433J3_126_901_n20, DP_OP_433J3_126_901_n15,
         DP_OP_433J3_126_901_n11, DP_OP_433J3_126_901_n7,
         DP_OP_433J3_126_901_n3, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n95, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n126, n127, n143, n146, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n884;
  wire   [2:0] StateMC;
  wire   [3:0] Debug_reg;
  wire   [8:0] Final_Exponent_reg;
  wire   [7:0] Op1_Mantissa_reg;
  wire   [7:0] Op2_Mantissa_reg;
  wire   [6:0] Final_Mantissa_reg;

  DFFRX1 T_reg_reg ( .D(n124), .CLK(CLK), .CLRB(n64), .Q(T_reg) );
  DFFRX1 exc_reg_reg_2_ ( .D(n667), .CLK(CLK), .CLRB(n64), .Q(n213), .QB(n74)
         );
  DFFRX1 StateMC_reg_0_ ( .D(n703), .CLK(CLK), .CLRB(n64), .Q(n66), .QB(
        StateMC[0]) );
  DFFRX1 StateMC_reg_1_ ( .D(N89), .CLK(CLK), .CLRB(n64), .Q(StateMC[1]), .QB(
        n57) );
  DFFRX1 StateMC_reg_2_ ( .D(N90), .CLK(CLK), .CLRB(n64), .Q(StateMC[2]), .QB(
        n65) );
  DFFRX1 Op1_Mantissa_reg_reg_0_ ( .D(n147), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[0]) );
  DFFRX1 Op1_Mantissa_reg_reg_1_ ( .D(n148), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[1]) );
  DFFRX1 Op1_Mantissa_reg_reg_2_ ( .D(n149), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[2]) );
  DFFRX1 Op1_Mantissa_reg_reg_3_ ( .D(n150), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[3]) );
  DFFRX1 Op1_Mantissa_reg_reg_4_ ( .D(n151), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[4]) );
  DFFRX1 Op1_Mantissa_reg_reg_5_ ( .D(n152), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[5]) );
  DFFRX1 Op1_Mantissa_reg_reg_6_ ( .D(n153), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[6]) );
  DFFRX1 Op1_Mantissa_reg_reg_7_ ( .D(n154), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[7]) );
  DFFRX1 Op2_Mantissa_reg_reg_0_ ( .D(n155), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[0]) );
  DFFRX1 Op2_Mantissa_reg_reg_1_ ( .D(n156), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[1]) );
  DFFRX1 Op2_Mantissa_reg_reg_2_ ( .D(n157), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[2]) );
  DFFRX1 Op2_Mantissa_reg_reg_3_ ( .D(n158), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[3]) );
  DFFRX1 Op2_Mantissa_reg_reg_4_ ( .D(n159), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[4]) );
  DFFRX1 Op2_Mantissa_reg_reg_5_ ( .D(n160), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[5]) );
  DFFRX1 Op2_Mantissa_reg_reg_6_ ( .D(n161), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[6]) );
  DFFRX1 Op2_Mantissa_reg_reg_7_ ( .D(n881), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[7]) );
  DFFRX1 exc_reg_reg_0_ ( .D(n882), .CLK(CLK), .CLRB(n64), .Q(n80), .QB(n215)
         );
  DFFRX1 Final_Exponent_reg_reg_8_ ( .D(n94), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[8]), .QB(n60) );
  DFFRX1 exc_reg_reg_1_ ( .D(n883), .CLK(CLK), .CLRB(n64), .Q(n77), .QB(n214)
         );
  DFFRX1 Final_Exponent_reg_reg_7_ ( .D(n872), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[7]), .QB(n72) );
  DFFRX1 Final_Exponent_reg_reg_6_ ( .D(n873), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[6]), .QB(n75) );
  DFFRX1 Final_Exponent_reg_reg_5_ ( .D(n874), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[5]), .QB(n69) );
  DFFRX1 Final_Exponent_reg_reg_4_ ( .D(n875), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[4]), .QB(n71) );
  DFFRX1 Final_Exponent_reg_reg_3_ ( .D(n876), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[3]), .QB(n59) );
  DFFRX1 Final_Exponent_reg_reg_2_ ( .D(n877), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[2]), .QB(n58) );
  DFFRX1 Final_Exponent_reg_reg_1_ ( .D(n878), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[1]), .QB(n61) );
  DFFRX1 Final_Exponent_reg_reg_0_ ( .D(n879), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[0]), .QB(n109) );
  DFFRX1 Debug_valid_reg_reg ( .D(n96), .CLK(CLK), .CLRB(n64), .Q(
        Debug_valid_reg) );
  DFFRX1 Final_Mantissa_reg_reg_0_ ( .D(n871), .CLK(CLK), .CLRB(n64), .Q(
        Final_Mantissa_reg[0]), .QB(n76) );
  DFFRX1 Final_Mantissa_reg_reg_1_ ( .D(n870), .CLK(CLK), .CLRB(n64), .Q(
        Final_Mantissa_reg[1]), .QB(n62) );
  DFFRX1 Final_Mantissa_reg_reg_2_ ( .D(n869), .CLK(CLK), .CLRB(n64), .Q(
        Final_Mantissa_reg[2]), .QB(n70) );
  DFFRX1 Final_Mantissa_reg_reg_3_ ( .D(n868), .CLK(CLK), .CLRB(n64), .Q(
        Final_Mantissa_reg[3]), .QB(n63) );
  DFFRX1 Final_Mantissa_reg_reg_4_ ( .D(n867), .CLK(CLK), .CLRB(n64), .Q(
        Final_Mantissa_reg[4]), .QB(n68) );
  DFFRX1 Final_Mantissa_reg_reg_5_ ( .D(n866), .CLK(CLK), .CLRB(n64), .Q(
        Final_Mantissa_reg[5]), .QB(n67) );
  DFFRX1 Final_Mantissa_reg_reg_6_ ( .D(n865), .CLK(CLK), .CLRB(n64), .Q(
        Final_Mantissa_reg[6]), .QB(n73) );
  DFFRX1 Final_Sign_reg_reg ( .D(n880), .CLK(CLK), .CLRB(n64), .Q(
        Final_Sign_reg), .QB(n78) );
  DFFRX1 G_reg_reg ( .D(n125), .CLK(CLK), .CLRB(n64), .Q(G_reg) );
  DFFRX1 Multi_datain1_reg_7_ ( .D(n163), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[7]) );
  DFFRX1 Multi_datain1_reg_6_ ( .D(n162), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[6]) );
  DFFRX1 Multi_datain1_reg_5_ ( .D(n133), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[5]) );
  DFFRX1 Multi_datain1_reg_4_ ( .D(n132), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[4]) );
  DFFRX1 Multi_datain1_reg_3_ ( .D(n131), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[3]) );
  DFFRX1 Multi_datain1_reg_2_ ( .D(n130), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[2]) );
  DFFRX1 Multi_datain1_reg_1_ ( .D(n129), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[1]) );
  DFFRX1 Multi_datain1_reg_0_ ( .D(n128), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[0]) );
  DFFRX1 Multi_datain2_reg_7_ ( .D(n141), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[7]) );
  DFFRX1 Multi_datain2_reg_6_ ( .D(n140), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[6]) );
  DFFRX1 Multi_datain2_reg_5_ ( .D(n139), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[5]) );
  DFFRX1 Multi_datain2_reg_4_ ( .D(n138), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[4]) );
  DFFRX1 Multi_datain2_reg_3_ ( .D(n137), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[3]) );
  DFFRX1 Multi_datain2_reg_2_ ( .D(n136), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[2]) );
  DFFRX1 Multi_datain2_reg_1_ ( .D(n135), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[1]) );
  DFFRX1 Multi_datain2_reg_0_ ( .D(n134), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[0]) );
  DFFRX1 Multi_valid_reg ( .D(n142), .CLK(CLK), .CLRB(n64), .QB(
        Multi_valid_BAR) );
  DFFRX1 ExcCheck_valid_reg ( .D(n864), .CLK(CLK), .CLRB(n64), .Q(
        ExcCheck_valid) );
  DFFRX1 Debug_reg_reg_3_ ( .D(n145), .CLK(CLK), .CLRB(n64), .Q(Debug_reg[3])
         );
  DFFRX1 Debug_reg_reg_2_ ( .D(n144), .CLK(CLK), .CLRB(n64), .Q(Debug_reg[2])
         );
  DFFRX1 Debug_reg_reg_1_ ( .D(n862), .CLK(CLK), .CLRB(n64), .Q(Debug_reg[1])
         );
  DFFRX1 Debug_reg_reg_0_ ( .D(n863), .CLK(CLK), .CLRB(n64), .Q(Debug_reg[0]), 
        .QB(n468) );
  NOR2X1 DP_OP_357J3_124_4634_U18 ( .IN1(Datain2[14]), .IN2(Datain1[14]), 
        .OUT(DP_OP_357J3_124_4634_n15) );
  NOR2X1 DP_OP_357J3_124_4634_U15 ( .IN1(Datain1[14]), .IN2(
        DP_OP_357J3_124_4634_n15), .OUT(DP_OP_357J3_124_4634_n13) );
  NOR2X1 DP_OP_357J3_124_4634_U14 ( .IN1(Datain2[14]), .IN2(
        DP_OP_357J3_124_4634_n15), .OUT(DP_OP_357J3_124_4634_n12) );
  NOR2X1 DP_OP_357J3_124_4634_U13 ( .IN1(DP_OP_357J3_124_4634_n13), .IN2(
        DP_OP_357J3_124_4634_n12), .OUT(DP_OP_357J3_124_4634_n17) );
  FULLADD DP_OP_357J3_124_4634_U12 ( .A(Datain1[7]), .B(Datain2[7]), .CIN(
        RSOP_428_C1_Z_0), .COUT(DP_OP_357J3_124_4634_n11), .SUM(N384) );
  FULLADD DP_OP_357J3_124_4634_U11 ( .A(DP_OP_357J3_124_4634_n11), .B(n146), 
        .CIN(DP_OP_357J3_124_4634_n29), .COUT(DP_OP_357J3_124_4634_n10), .SUM(
        N385) );
  FULLADD DP_OP_357J3_124_4634_U10 ( .A(DP_OP_357J3_124_4634_n27), .B(
        DP_OP_357J3_124_4634_n28), .CIN(DP_OP_357J3_124_4634_n10), .COUT(
        DP_OP_357J3_124_4634_n9), .SUM(N386) );
  FULLADD DP_OP_357J3_124_4634_U9 ( .A(DP_OP_357J3_124_4634_n25), .B(
        DP_OP_357J3_124_4634_n26), .CIN(DP_OP_357J3_124_4634_n9), .COUT(
        DP_OP_357J3_124_4634_n8), .SUM(N387) );
  FULLADD DP_OP_357J3_124_4634_U8 ( .A(DP_OP_357J3_124_4634_n23), .B(
        DP_OP_357J3_124_4634_n24), .CIN(DP_OP_357J3_124_4634_n8), .COUT(
        DP_OP_357J3_124_4634_n7), .SUM(N388) );
  FULLADD DP_OP_357J3_124_4634_U7 ( .A(DP_OP_357J3_124_4634_n21), .B(
        DP_OP_357J3_124_4634_n22), .CIN(DP_OP_357J3_124_4634_n7), .COUT(
        DP_OP_357J3_124_4634_n6), .SUM(N389) );
  FULLADD DP_OP_357J3_124_4634_U6 ( .A(DP_OP_357J3_124_4634_n19), .B(
        DP_OP_357J3_124_4634_n20), .CIN(DP_OP_357J3_124_4634_n6), .COUT(
        DP_OP_357J3_124_4634_n5), .SUM(N390) );
  FULLADD DP_OP_357J3_124_4634_U5 ( .A(DP_OP_357J3_124_4634_n18), .B(
        DP_OP_357J3_124_4634_n17), .CIN(DP_OP_357J3_124_4634_n5), .COUT(
        DP_OP_357J3_124_4634_n4), .SUM(N391) );
  NOR2X1 DP_OP_357J3_124_4634_U4 ( .IN1(DP_OP_357J3_124_4634_n4), .IN2(n123), 
        .OUT(DP_OP_357J3_124_4634_n3) );
  NOR2X1 DP_OP_357J3_124_4634_U3 ( .IN1(DP_OP_357J3_124_4634_n4), .IN2(
        DP_OP_357J3_124_4634_n3), .OUT(DP_OP_357J3_124_4634_n2) );
  NOR2X1 DP_OP_357J3_124_4634_U2 ( .IN1(n123), .IN2(DP_OP_357J3_124_4634_n3), 
        .OUT(DP_OP_357J3_124_4634_n1) );
  NOR2X1 DP_OP_357J3_124_4634_U1 ( .IN1(DP_OP_357J3_124_4634_n2), .IN2(
        DP_OP_357J3_124_4634_n1), .OUT(N392) );
  NOR2X1 DP_OP_433J3_126_901_U34 ( .IN1(n119), .IN2(DP_OP_433J3_126_901_n23), 
        .OUT(DP_OP_433J3_126_901_n21) );
  NOR2X1 DP_OP_433J3_126_901_U33 ( .IN1(Final_Exponent_reg[0]), .IN2(
        DP_OP_433J3_126_901_n23), .OUT(DP_OP_433J3_126_901_n20) );
  NOR2X1 DP_OP_433J3_126_901_U32 ( .IN1(DP_OP_433J3_126_901_n21), .IN2(
        DP_OP_433J3_126_901_n20), .OUT(C276_DATA3_0) );
  FULLADD DP_OP_433J3_126_901_U31 ( .A(n118), .B(n116), .CIN(n108), .COUT(
        DP_OP_433J3_126_901_n30), .SUM(C276_DATA3_1) );
  FULLADD DP_OP_433J3_126_901_U30 ( .A(n302), .B(Final_Exponent_reg[2]), .CIN(
        n106), .COUT(DP_OP_433J3_126_901_n29), .SUM(C276_DATA3_2) );
  FULLADD DP_OP_433J3_126_901_U29 ( .A(n117), .B(Final_Exponent_reg[3]), .CIN(
        n107), .COUT(DP_OP_433J3_126_901_n28), .SUM(C276_DATA3_3) );
  NOR2X1 DP_OP_433J3_126_901_U16 ( .IN1(Final_Exponent_reg[6]), .IN2(n111), 
        .OUT(DP_OP_433J3_126_901_n11) );
  NOR2X1 DP_OP_433J3_126_901_U10 ( .IN1(Final_Exponent_reg[7]), .IN2(n121), 
        .OUT(DP_OP_433J3_126_901_n7) );
  NOR2X1 DP_OP_433J3_126_901_U4 ( .IN1(n122), .IN2(Final_Exponent_reg[8]), 
        .OUT(DP_OP_433J3_126_901_n3) );
  BUF4X U3 ( .IN(DP_OP_433J3_126_901_n29), .OUT(n107) );
  BUF4X U4 ( .IN(DP_OP_433J3_126_901_n30), .OUT(n106) );
  AOI21 U5 ( .IN1(Final_Exponent_reg[4]), .IN2(DP_OP_433J3_126_901_n28), .IN3(
        n56), .OUT(n1) );
  NAND3X1 U6 ( .IN1(n270), .IN2(n269), .IN3(n283), .OUT(n2) );
  AOI21 U7 ( .IN1(n500), .IN2(N388), .IN3(n2), .OUT(n3) );
  OAI21 U8 ( .IN1(n4), .IN2(n1), .IN3(n3), .OUT(n5) );
  AOI21 U9 ( .IN1(n496), .IN2(Final_Exponent_reg[4]), .IN3(n287), .OUT(n6) );
  OAI21 U10 ( .IN1(n126), .IN2(n7), .IN3(n6), .OUT(n875) );
  INVX1 U11 ( .IN(n339), .OUT(n4) );
  INVX1 U12 ( .IN(n5), .OUT(n7) );
  INVX1 U13 ( .IN(n393), .OUT(n8) );
  NAND3X1 U14 ( .IN1(n392), .IN2(n650), .IN3(n394), .OUT(n9) );
  NOR2X1 U15 ( .IN1(n8), .IN2(n9), .OUT(n10) );
  NOR2X1 U16 ( .IN1(n409), .IN2(n387), .OUT(n11) );
  NAND3X1 U17 ( .IN1(n389), .IN2(n388), .IN3(n11), .OUT(n12) );
  NAND2X1 U18 ( .IN1(n390), .IN2(n391), .OUT(n13) );
  NAND3X1 U19 ( .IN1(n448), .IN2(n449), .IN3(n13), .OUT(n14) );
  OAI21 U20 ( .IN1(n12), .IN2(n14), .IN3(n55), .OUT(n15) );
  NAND3X1 U21 ( .IN1(n395), .IN2(n10), .IN3(n15), .OUT(n402) );
  INVX1 U22 ( .IN(n339), .OUT(n16) );
  AOI21 U23 ( .IN1(Final_Exponent_reg[5]), .IN2(n120), .IN3(
        DP_OP_433J3_126_901_n15), .OUT(n17) );
  AOI21 U24 ( .IN1(N389), .IN2(n500), .IN3(n277), .OUT(n18) );
  OAI21 U25 ( .IN1(n16), .IN2(n17), .IN3(n18), .OUT(n19) );
  INVX1 U26 ( .IN(n19), .OUT(n20) );
  AOI21 U27 ( .IN1(n293), .IN2(Final_Exponent_reg[5]), .IN3(n340), .OUT(n21)
         );
  OAI21 U28 ( .IN1(n126), .IN2(n20), .IN3(n21), .OUT(n874) );
  NAND3X1 U29 ( .IN1(n446), .IN2(n441), .IN3(n448), .OUT(n464) );
  AOI21 U30 ( .IN1(n111), .IN2(Final_Exponent_reg[6]), .IN3(
        DP_OP_433J3_126_901_n11), .OUT(n22) );
  INVX1 U31 ( .IN(n339), .OUT(n23) );
  AOI21 U32 ( .IN1(n286), .IN2(Final_Exponent_reg[6]), .IN3(n285), .OUT(n24)
         );
  OAI21 U33 ( .IN1(n22), .IN2(n23), .IN3(n24), .OUT(n25) );
  AOI21 U34 ( .IN1(n500), .IN2(N390), .IN3(n25), .OUT(n26) );
  AOI21 U35 ( .IN1(n496), .IN2(Final_Exponent_reg[6]), .IN3(n287), .OUT(n27)
         );
  OAI21 U36 ( .IN1(n126), .IN2(n26), .IN3(n27), .OUT(n873) );
  AOI21 U37 ( .IN1(n122), .IN2(Final_Exponent_reg[8]), .IN3(
        DP_OP_433J3_126_901_n3), .OUT(n28) );
  INVX1 U38 ( .IN(n28), .OUT(C276_DATA3_8) );
  NAND3X1 U39 ( .IN1(n66), .IN2(n65), .IN3(StateMC[1]), .OUT(n777) );
  NAND3X1 U40 ( .IN1(n378), .IN2(n406), .IN3(n388), .OUT(n29) );
  AOI21 U41 ( .IN1(n427), .IN2(n379), .IN3(n29), .OUT(n30) );
  AOI21 U42 ( .IN1(n405), .IN2(n383), .IN3(n391), .OUT(n31) );
  NAND3X1 U43 ( .IN1(n30), .IN2(n384), .IN3(n31), .OUT(n32) );
  AOI21 U44 ( .IN1(n116), .IN2(n32), .IN3(C1_Z_1), .OUT(n752) );
  NAND3X1 U45 ( .IN1(Final_Exponent_reg[6]), .IN2(Final_Exponent_reg[5]), 
        .IN3(n272), .OUT(n281) );
  NAND3X1 U46 ( .IN1(n214), .IN2(n215), .IN3(n213), .OUT(n789) );
  AOI22 U47 ( .IN1(Datain1[5]), .IN2(n497), .IN3(Datain2[5]), .IN4(n498), 
        .OUT(n33) );
  AOI22 U48 ( .IN1(n745), .IN2(Multi_dataout[13]), .IN3(n744), .IN4(
        Multi_dataout[12]), .OUT(n34) );
  INVX1 U49 ( .IN(n740), .OUT(n35) );
  AOI21 U50 ( .IN1(Final_Mantissa_reg[5]), .IN2(n35), .IN3(n512), .OUT(n36) );
  OAI21 U51 ( .IN1(Final_Mantissa_reg[5]), .IN2(n35), .IN3(n36), .OUT(n37) );
  NAND3X1 U52 ( .IN1(n33), .IN2(n34), .IN3(n37), .OUT(n38) );
  INVX1 U53 ( .IN(n400), .OUT(n39) );
  AOI22 U54 ( .IN1(n400), .IN2(n742), .IN3(n741), .IN4(n39), .OUT(n40) );
  AOI22 U55 ( .IN1(n114), .IN2(Multi_dataout[9]), .IN3(n113), .IN4(
        Multi_dataout[10]), .OUT(n41) );
  OAI21 U56 ( .IN1(n509), .IN2(n760), .IN3(n41), .OUT(n42) );
  AOI22 U57 ( .IN1(n743), .IN2(n762), .IN3(n764), .IN4(n42), .OUT(n43) );
  OAI21 U58 ( .IN1(n766), .IN2(n40), .IN3(n43), .OUT(n44) );
  OAI21 U59 ( .IN1(n38), .IN2(n44), .IN3(RSTn), .OUT(n45) );
  OAI21 U60 ( .IN1(n771), .IN2(n67), .IN3(n45), .OUT(n866) );
  AOI21 U61 ( .IN1(Final_Exponent_reg[7]), .IN2(n121), .IN3(
        DP_OP_433J3_126_901_n7), .OUT(n46) );
  AOI21 U62 ( .IN1(N391), .IN2(n500), .IN3(n292), .OUT(n47) );
  OAI21 U63 ( .IN1(n48), .IN2(n46), .IN3(n47), .OUT(n49) );
  AOI21 U64 ( .IN1(n293), .IN2(Final_Exponent_reg[7]), .IN3(n340), .OUT(n50)
         );
  OAI21 U65 ( .IN1(n126), .IN2(n51), .IN3(n50), .OUT(n872) );
  INVX1 U66 ( .IN(n339), .OUT(n48) );
  INVX1 U67 ( .IN(n49), .OUT(n51) );
  INVX4 U68 ( .IN(Exc_Ack_BAR), .OUT(n52) );
  INVX1 U69 ( .IN(Multi_dataout[13]), .OUT(n455) );
  INVX1 U70 ( .IN(n329), .OUT(n94) );
  INVX1 U71 ( .IN(n478), .OUT(n863) );
  NANDX2 U72 ( .IN1(n250), .IN2(n266), .OUT(n879) );
  NAND2X1 U73 ( .IN1(n702), .IN2(n701), .OUT(n705) );
  NAND2X1 U74 ( .IN1(n339), .IN2(C276_DATA3_2), .OUT(n262) );
  INVX1 U75 ( .IN(n825), .OUT(n145) );
  NANDX2 U76 ( .IN1(n782), .IN2(n486), .OUT(n766) );
  INVX1 U77 ( .IN(n471), .OUT(n472) );
  NANDX2 U78 ( .IN1(n495), .IN2(n651), .OUT(n782) );
  INVX1 U79 ( .IN(n351), .OUT(n651) );
  NAND2X1 U80 ( .IN1(n317), .IN2(n316), .OUT(n318) );
  INVX1 U81 ( .IN(n375), .OUT(n376) );
  INVX1 U82 ( .IN(n419), .OUT(n423) );
  NAND2X1 U83 ( .IN1(n315), .IN2(n433), .OUT(n316) );
  INVX1 U84 ( .IN(n232), .OUT(n233) );
  NANDX2 U85 ( .IN1(n303), .IN2(n207), .OUT(n372) );
  INVX1 U86 ( .IN(n453), .OUT(n462) );
  INVX1 U87 ( .IN(n303), .OUT(n494) );
  NAND2X1 U88 ( .IN1(n392), .IN2(n303), .OUT(n308) );
  NAND2X1 U89 ( .IN1(n362), .IN2(n361), .OUT(n364) );
  INVX1 U90 ( .IN(n439), .OUT(n440) );
  NAND2X1 U91 ( .IN1(n465), .IN2(n432), .OUT(n457) );
  INVX1 U92 ( .IN(n582), .OUT(n587) );
  NAND2X1 U93 ( .IN1(n474), .IN2(n486), .OUT(n404) );
  NAND2X1 U94 ( .IN1(n500), .IN2(N387), .OUT(n336) );
  NANDX2 U95 ( .IN1(n311), .IN2(n299), .OUT(n206) );
  INVX1 U96 ( .IN(n841), .OUT(n137) );
  NANDX2 U97 ( .IN1(n368), .IN2(n365), .OUT(n393) );
  INVX1 U98 ( .IN(n839), .OUT(n139) );
  INVX1 U99 ( .IN(n843), .OUT(n135) );
  INVX1 U100 ( .IN(n849), .OUT(n129) );
  INVX1 U101 ( .IN(n837), .OUT(n141) );
  INVX1 U102 ( .IN(n838), .OUT(n140) );
  INVX1 U103 ( .IN(n847), .OUT(n131) );
  INVX1 U104 ( .IN(n844), .OUT(n134) );
  INVX1 U105 ( .IN(n840), .OUT(n138) );
  INVX1 U106 ( .IN(n852), .OUT(n128) );
  INVX1 U107 ( .IN(n848), .OUT(n130) );
  INVX1 U108 ( .IN(n842), .OUT(n136) );
  INVX1 U109 ( .IN(n273), .OUT(n647) );
  INVX1 U110 ( .IN(n492), .OUT(n628) );
  INVX1 U111 ( .IN(n846), .OUT(n132) );
  INVX1 U112 ( .IN(n845), .OUT(n133) );
  INVX1 U113 ( .IN(n459), .OUT(n355) );
  NAND2X1 U114 ( .IN1(n500), .IN2(N384), .OUT(n243) );
  INVX1 U115 ( .IN(n454), .OUT(n179) );
  INVX1 U116 ( .IN(n804), .OUT(n162) );
  INVX1 U117 ( .IN(n801), .OUT(n163) );
  NAND2X1 U118 ( .IN1(n354), .IN2(n353), .OUT(n459) );
  NANDX2 U119 ( .IN1(Final_Exponent_reg[7]), .IN2(n289), .OUT(n288) );
  NAND2X1 U120 ( .IN1(n596), .IN2(n595), .OUT(n597) );
  NAND2X1 U121 ( .IN1(n484), .IN2(n483), .OUT(n485) );
  INVX1 U122 ( .IN(n346), .OUT(n347) );
  NAND2X1 U123 ( .IN1(n669), .IN2(n746), .OUT(n861) );
  INVX1 U124 ( .IN(n621), .OUT(n881) );
  NAND2X1 U125 ( .IN1(n503), .IN2(n821), .OUT(n659) );
  NAND2X1 U126 ( .IN1(n452), .IN2(n489), .OUT(n477) );
  INVX1 U127 ( .IN(n816), .OUT(n150) );
  INVX1 U128 ( .IN(n815), .OUT(n151) );
  INVX1 U129 ( .IN(n817), .OUT(n149) );
  INVX1 U130 ( .IN(n814), .OUT(n152) );
  INVX1 U131 ( .IN(n818), .OUT(n148) );
  INVX1 U132 ( .IN(n820), .OUT(n147) );
  INVX1 U133 ( .IN(n813), .OUT(n153) );
  INVX1 U134 ( .IN(n812), .OUT(n154) );
  INVX1 U135 ( .IN(n811), .OUT(n155) );
  INVX1 U136 ( .IN(n810), .OUT(n156) );
  INVX1 U137 ( .IN(n809), .OUT(n157) );
  NAND2X1 U138 ( .IN1(n504), .IN2(n610), .OUT(n346) );
  INVX1 U139 ( .IN(n808), .OUT(n158) );
  NANDX2 U140 ( .IN1(n61), .IN2(n360), .OUT(n356) );
  INVX1 U141 ( .IN(n807), .OUT(n159) );
  INVX1 U142 ( .IN(n806), .OUT(n160) );
  INVX1 U143 ( .IN(n805), .OUT(n161) );
  INVX1 U144 ( .IN(n610), .OUT(n168) );
  INVX1 U145 ( .IN(n354), .OUT(n190) );
  NAND2X1 U146 ( .IN1(n639), .IN2(n709), .OUT(n746) );
  NAND2X1 U147 ( .IN1(Multi_dataout[14]), .IN2(n507), .OUT(n781) );
  INVX4 U148 ( .IN(Multi_dataout[1]), .OUT(n225) );
  NANDX2 U149 ( .IN1(Multi_dataout[4]), .IN2(n212), .OUT(n200) );
  INVX1 U150 ( .IN(n799), .OUT(n800) );
  INVX1 U151 ( .IN(n553), .OUT(n557) );
  INVX1 U152 ( .IN(Multi_dataout[14]), .OUT(n317) );
  INVX1 U153 ( .IN(n484), .OUT(n422) );
  NAND2X1 U154 ( .IN1(n854), .IN2(n853), .OUT(n627) );
  NANDX2 U155 ( .IN1(n646), .IN2(Final_Exponent_reg[4]), .OUT(n278) );
  NANDX2 U156 ( .IN1(n58), .IN2(n366), .OUT(n368) );
  NAND2X1 U157 ( .IN1(n631), .IN2(n511), .OUT(n602) );
  INVX1 U158 ( .IN(n633), .OUT(n238) );
  NAND2X1 U159 ( .IN1(n634), .IN2(n240), .OUT(n333) );
  NAND2X1 U160 ( .IN1(n728), .IN2(Final_Mantissa_reg[4]), .OUT(n740) );
  NAND2X1 U161 ( .IN1(n52), .IN2(n630), .OUT(n548) );
  INVX1 U162 ( .IN(Exc[2]), .OUT(n590) );
  NAND2X1 U163 ( .IN1(n779), .IN2(n581), .OUT(n584) );
  INVX1 U164 ( .IN(n634), .OUT(n630) );
  NANDX2 U165 ( .IN1(n59), .IN2(n227), .OUT(n358) );
  INVX1 U166 ( .IN(n629), .OUT(n240) );
  INVX1 U167 ( .IN(n559), .OUT(Debug[1]) );
  INVX1 U168 ( .IN(n479), .OUT(Debug[0]) );
  INVX1 U169 ( .IN(n561), .OUT(Debug[3]) );
  INVX1 U170 ( .IN(n564), .OUT(Debug[4]) );
  INVX1 U171 ( .IN(n560), .OUT(Debug[2]) );
  INVX4 U172 ( .IN(n581), .OUT(n53) );
  INVX1 U173 ( .IN(n642), .OUT(n186) );
  NAND2X1 U174 ( .IN1(n583), .IN2(n543), .OUT(n544) );
  NANDX2 U175 ( .IN1(n693), .IN2(Final_Mantissa_reg[2]), .OUT(n707) );
  NANDX2 U176 ( .IN1(n166), .IN2(StateMC[0]), .OUT(n585) );
  INVX1 U177 ( .IN(n778), .OUT(n170) );
  INVX1 U178 ( .IN(n52), .OUT(n543) );
  INVX1 U179 ( .IN(DP_OP_357J3_124_4634_n15), .OUT(n123) );
  INVX1 U180 ( .IN(n772), .OUT(n166) );
  INVX4 U181 ( .IN(Datain2[7]), .OUT(n523) );
  NAND2X1 U182 ( .IN1(n481), .IN2(n420), .OUT(n563) );
  INVX1 U183 ( .IN(n420), .OUT(n421) );
  INVX1 U184 ( .IN(Datain1[9]), .OUT(n529) );
  NANDX2 U185 ( .IN1(StateMC[2]), .IN2(StateMC[1]), .OUT(n171) );
  INVX1 U186 ( .IN(Datain2[10]), .OUT(n520) );
  INVX1 U187 ( .IN(Datain2[11]), .OUT(n521) );
  NANDX2 U188 ( .IN1(Datain1[11]), .IN2(Datain2[11]), .OUT(n92) );
  NANDX2 U189 ( .IN1(Datain1[10]), .IN2(Datain2[10]), .OUT(n88) );
  NANDX2 U190 ( .IN1(n57), .IN2(n65), .OUT(n772) );
  INVX1 U191 ( .IN(n58), .OUT(n55) );
  INVX1 U192 ( .IN(Datain1[8]), .OUT(n530) );
  INVX1 U193 ( .IN(Datain2[8]), .OUT(n524) );
  INVX1 U194 ( .IN(Datain1[11]), .OUT(n533) );
  INVX1 U195 ( .IN(Datain1[12]), .OUT(n532) );
  NANDX2 U196 ( .IN1(n61), .IN2(n109), .OUT(n195) );
  NANDX2 U197 ( .IN1(Mode[0]), .IN2(Mode[2]), .OUT(n481) );
  NANDX2 U198 ( .IN1(StateMC[0]), .IN2(n505), .OUT(n604) );
  NANDX2 U199 ( .IN1(n66), .IN2(n505), .OUT(n581) );
  NOR2X1 U200 ( .IN1(Final_Exponent_reg[4]), .IN2(DP_OP_433J3_126_901_n28), 
        .OUT(n56) );
  INVX1 U201 ( .IN(n56), .OUT(n120) );
  INVX1 U202 ( .IN(n441), .OUT(n391) );
  NAND2X1 U203 ( .IN1(RSTn), .IN2(n836), .OUT(n833) );
  NAND2X1 U204 ( .IN1(n831), .IN2(n830), .OUT(n144) );
  INVX1 U205 ( .IN(n771), .OUT(n704) );
  NAND2X1 U206 ( .IN1(RSTn), .IN2(n772), .OUT(n853) );
  INVX1 U207 ( .IN(n746), .OUT(n747) );
  INVX1 U208 ( .IN(Multi_dataout[0]), .OUT(n755) );
  NANDX2 U209 ( .IN1(n257), .IN2(n266), .OUT(n878) );
  NAND2X1 U210 ( .IN1(n339), .IN2(C276_DATA3_1), .OUT(n254) );
  NAND2X1 U211 ( .IN1(n647), .IN2(n646), .OUT(n648) );
  NANDX2 U212 ( .IN1(n298), .IN2(n373), .OUT(n235) );
  NANDX2 U213 ( .IN1(n116), .IN2(Final_Exponent_reg[0]), .OUT(n642) );
  NANDX2 U214 ( .IN1(n748), .IN2(Final_Mantissa_reg[6]), .OUT(n639) );
  NAND2X1 U215 ( .IN1(n171), .IN2(n170), .OUT(n172) );
  INVX1 U216 ( .IN(n268), .OUT(n269) );
  INVX4 U217 ( .IN(n294), .OUT(n350) );
  NAND2X1 U218 ( .IN1(n442), .IN2(n449), .OUT(n460) );
  NANDX2 U219 ( .IN1(RSTn), .IN2(n172), .OUT(n884) );
  NANDX2 U220 ( .IN1(RSTn), .IN2(n503), .OUT(n854) );
  INVX4 U221 ( .IN(Multi_dataout[15]), .OUT(n507) );
  NANDX2 U222 ( .IN1(n370), .IN2(n384), .OUT(n371) );
  NANDX2 U223 ( .IN1(n255), .IN2(n254), .OUT(n256) );
  NANDX2 U224 ( .IN1(n199), .IN2(n227), .OUT(n209) );
  INVX4 U225 ( .IN(n854), .OUT(n319) );
  NANDX2 U226 ( .IN1(n164), .IN2(n346), .OUT(n165) );
  NAND2X1 U227 ( .IN1(Datain1[8]), .IN2(Datain2[8]), .OUT(n81) );
  NANDX2 U228 ( .IN1(n412), .IN2(n406), .OUT(n314) );
  NANDX2 U229 ( .IN1(Multi_dataout[5]), .IN2(n482), .OUT(n412) );
  NANDX2 U230 ( .IN1(n319), .IN2(n836), .OUT(n452) );
  INVX4 U231 ( .IN(n766), .OUT(n399) );
  NANDX2 U232 ( .IN1(n263), .IN2(n262), .OUT(n264) );
  NANDX2 U233 ( .IN1(n421), .IN2(n504), .OUT(n484) );
  NANDX2 U234 ( .IN1(n180), .IN2(n366), .OUT(n185) );
  NAND2X1 U235 ( .IN1(Final_Exponent_reg[2]), .IN2(n186), .OUT(n644) );
  NAND2X1 U236 ( .IN1(Datain1[9]), .IN2(Datain2[9]), .OUT(n84) );
  NAND2X1 U237 ( .IN1(Datain1[12]), .IN2(Datain2[12]), .OUT(n97) );
  INVX4 U238 ( .IN(n709), .OUT(n512) );
  NANDX2 U239 ( .IN1(n350), .IN2(n373), .OUT(n295) );
  NANDX2 U240 ( .IN1(n507), .IN2(n317), .OUT(n169) );
  NAND2X1 U241 ( .IN1(n344), .IN2(n776), .OUT(n321) );
  NANDX2 U242 ( .IN1(n201), .IN2(n386), .OUT(n202) );
  BUF4X U243 ( .IN(n819), .OUT(n112) );
  BUF4X U244 ( .IN(n851), .OUT(n115) );
  INVX4 U245 ( .IN(n612), .OUT(n598) );
  INVX4 U246 ( .IN(n349), .OUT(n491) );
  INVX4 U247 ( .IN(n618), .OUT(n127) );
  NAND2X1 U248 ( .IN1(Datain1[13]), .IN2(Datain2[13]), .OUT(n101) );
  INVX4 U249 ( .IN(n295), .OUT(n296) );
  NANDX2 U250 ( .IN1(n507), .IN2(n318), .OUT(n776) );
  INVX4 U251 ( .IN(n202), .OUT(n203) );
  NANDX2 U252 ( .IN1(n465), .IN2(n434), .OUT(n480) );
  NANDX2 U253 ( .IN1(n726), .IN2(n788), .OUT(n711) );
  NANDX2 U254 ( .IN1(RSTn), .IN2(n248), .OUT(n271) );
  NANDX2 U255 ( .IN1(n821), .IN2(n776), .OUT(n640) );
  NANDX2 U256 ( .IN1(n69), .IN2(n56), .OUT(n111) );
  NANDX2 U257 ( .IN1(n109), .IN2(C1_Z_0), .OUT(n108) );
  NANDX2 U258 ( .IN1(n296), .IN2(n395), .OUT(n297) );
  NANDX2 U259 ( .IN1(n219), .IN2(n304), .OUT(n220) );
  NANDX2 U260 ( .IN1(n193), .IN2(n306), .OUT(n194) );
  INVX1 U261 ( .IN(n430), .OUT(n380) );
  INVX4 U262 ( .IN(n368), .OUT(n360) );
  NANDX2 U263 ( .IN1(n482), .IN2(n446), .OUT(n222) );
  INVX4 U264 ( .IN(n200), .OUT(n205) );
  INVX4 U265 ( .IN(n216), .OUT(n217) );
  NANDX2 U266 ( .IN1(n430), .IN2(n203), .OUT(n204) );
  INVX4 U267 ( .IN(Multi_dataout[10]), .OUT(n176) );
  NANDX2 U268 ( .IN1(n344), .IN2(Multi_dataout[15]), .OUT(n167) );
  INVX4 U269 ( .IN(n436), .OUT(n823) );
  NANDX2 U270 ( .IN1(n662), .IN2(n661), .OUT(n733) );
  NANDX2 U271 ( .IN1(n654), .IN2(n653), .OUT(n725) );
  NANDX2 U272 ( .IN1(n726), .IN2(n741), .OUT(n684) );
  INVX4 U273 ( .IN(n698), .OUT(n726) );
  NANDX2 U274 ( .IN1(n399), .IN2(n400), .OUT(n698) );
  NANDX2 U275 ( .IN1(n677), .IN2(n676), .OUT(n678) );
  NANDX2 U276 ( .IN1(n690), .IN2(n689), .OUT(n761) );
  NANDX2 U277 ( .IN1(n680), .IN2(n679), .OUT(n743) );
  INVX4 U278 ( .IN(n398), .OUT(n762) );
  NANDX2 U279 ( .IN1(n682), .IN2(n681), .OUT(n742) );
  INVX4 U280 ( .IN(n396), .OUT(n764) );
  NANDX2 U281 ( .IN1(n785), .IN2(n784), .OUT(n857) );
  INVX4 U282 ( .IN(n402), .OUT(n400) );
  NANDX2 U283 ( .IN1(n692), .IN2(n691), .OUT(n756) );
  NANDX2 U284 ( .IN1(n793), .IN2(n792), .OUT(n855) );
  NANDX2 U285 ( .IN1(n719), .IN2(n718), .OUT(n787) );
  INVX4 U286 ( .IN(n683), .OUT(n717) );
  NANDX2 U287 ( .IN1(n652), .IN2(n752), .OUT(n683) );
  INVX4 U288 ( .IN(n754), .OUT(n652) );
  INVX4 U289 ( .IN(n760), .OUT(n716) );
  NANDX2 U290 ( .IN1(n754), .IN2(n752), .OUT(n760) );
  NANDX2 U291 ( .IN1(n377), .IN2(n376), .OUT(n754) );
  NANDX2 U292 ( .IN1(n490), .IN2(n469), .OUT(n483) );
  INVX4 U293 ( .IN(n171), .OUT(n505) );
  NANDX2 U294 ( .IN1(n266), .IN2(n265), .OUT(n877) );
  INVX4 U295 ( .IN(n333), .OUT(n497) );
  NANDX2 U296 ( .IN1(n249), .IN2(n271), .OUT(n340) );
  NANDX2 U297 ( .IN1(n655), .IN2(n345), .OUT(n248) );
  NANDX2 U298 ( .IN1(n589), .IN2(n511), .OUT(n655) );
  NAND2X1 U299 ( .IN1(RSTn), .IN2(n267), .OUT(n249) );
  INVX4 U300 ( .IN(n884), .OUT(n496) );
  INVX4 U301 ( .IN(n239), .OUT(n498) );
  NANDX2 U302 ( .IN1(n238), .IN2(n511), .OUT(n239) );
  NANDX2 U303 ( .IN1(n583), .IN2(n52), .OUT(n632) );
  NANDX2 U304 ( .IN1(n579), .IN2(n52), .OUT(n629) );
  INVX4 U305 ( .IN(n668), .OUT(n821) );
  NANDX2 U306 ( .IN1(n344), .IN2(Multi_ack), .OUT(n668) );
  INVX4 U307 ( .IN(n279), .OUT(n649) );
  NANDX2 U308 ( .IN1(n660), .IN2(n241), .OUT(n279) );
  NANDX2 U309 ( .IN1(n469), .IN2(n502), .OUT(n660) );
  NANDX2 U310 ( .IN1(n486), .IN2(n322), .OUT(n237) );
  NANDX2 U311 ( .IN1(n469), .IN2(n323), .OUT(n385) );
  INVX4 U312 ( .IN(n794), .OUT(n469) );
  NANDX2 U313 ( .IN1(n428), .IN2(n445), .OUT(n453) );
  INVX4 U314 ( .IN(n474), .OUT(n490) );
  NANDX2 U315 ( .IN1(n403), .IN2(n465), .OUT(n474) );
  INVX4 U316 ( .IN(RSTn), .OUT(n126) );
  NANDX2 U317 ( .IN1(n82), .IN2(n83), .OUT(DP_OP_357J3_124_4634_n29) );
  INVX4 U318 ( .IN(n146), .OUT(RSOP_428_C1_Z_0) );
  NANDX2 U319 ( .IN1(n143), .IN2(n127), .OUT(n146) );
  INVX4 U320 ( .IN(n81), .OUT(DP_OP_357J3_124_4634_n28) );
  NANDX2 U321 ( .IN1(n86), .IN2(n87), .OUT(DP_OP_357J3_124_4634_n27) );
  INVX4 U322 ( .IN(n84), .OUT(DP_OP_357J3_124_4634_n26) );
  NANDX2 U323 ( .IN1(n90), .IN2(n91), .OUT(DP_OP_357J3_124_4634_n25) );
  INVX4 U324 ( .IN(n88), .OUT(DP_OP_357J3_124_4634_n24) );
  NANDX2 U325 ( .IN1(n93), .IN2(n95), .OUT(DP_OP_357J3_124_4634_n23) );
  INVX4 U326 ( .IN(n92), .OUT(DP_OP_357J3_124_4634_n22) );
  NANDX2 U327 ( .IN1(n99), .IN2(n100), .OUT(DP_OP_357J3_124_4634_n21) );
  INVX4 U328 ( .IN(n97), .OUT(DP_OP_357J3_124_4634_n20) );
  NANDX2 U329 ( .IN1(n104), .IN2(n105), .OUT(DP_OP_357J3_124_4634_n19) );
  INVX4 U330 ( .IN(n101), .OUT(DP_OP_357J3_124_4634_n18) );
  NANDX2 U331 ( .IN1(n504), .IN2(n168), .OUT(n596) );
  INVX4 U332 ( .IN(n473), .OUT(n326) );
  NANDX2 U333 ( .IN1(n325), .IN2(n324), .OUT(n473) );
  INVX4 U334 ( .IN(C1_Z_1), .OUT(n118) );
  NANDX2 U335 ( .IN1(n309), .IN2(n373), .OUT(C1_Z_1) );
  INVX4 U336 ( .IN(n299), .OUT(n493) );
  INVX4 U337 ( .IN(C1_Z_3), .OUT(n117) );
  INVX4 U338 ( .IN(n297), .OUT(n310) );
  NANDX2 U339 ( .IN1(n236), .IN2(n495), .OUT(n322) );
  NANDX2 U340 ( .IN1(n394), .IN2(n395), .OUT(n300) );
  NANDX2 U341 ( .IN1(n234), .IN2(n405), .OUT(n395) );
  INVX4 U342 ( .IN(n448), .OUT(n405) );
  INVX4 U343 ( .IN(n383), .OUT(n234) );
  NANDX2 U344 ( .IN1(n230), .IN2(n229), .OUT(n383) );
  NANDX2 U345 ( .IN1(n228), .IN2(n227), .OUT(n230) );
  NANDX2 U346 ( .IN1(n229), .IN2(n415), .OUT(n394) );
  INVX4 U347 ( .IN(n449), .OUT(n415) );
  INVX4 U348 ( .IN(n390), .OUT(n229) );
  NANDX2 U349 ( .IN1(n223), .IN2(n391), .OUT(n373) );
  NANDX2 U350 ( .IN1(n221), .IN2(n358), .OUT(n390) );
  INVX4 U351 ( .IN(n220), .OUT(n298) );
  NANDX2 U352 ( .IN1(n363), .IN2(n218), .OUT(n304) );
  INVX4 U353 ( .IN(n210), .OUT(n363) );
  NANDX2 U354 ( .IN1(n198), .IN2(n427), .OUT(n299) );
  INVX4 U355 ( .IN(n379), .OUT(n198) );
  NANDX2 U356 ( .IN1(n196), .IN2(n368), .OUT(n379) );
  NANDX2 U357 ( .IN1(n228), .IN2(n366), .OUT(n196) );
  INVX4 U358 ( .IN(n195), .OUT(n228) );
  INVX4 U359 ( .IN(n194), .OUT(n311) );
  NANDX2 U360 ( .IN1(n192), .IN2(n352), .OUT(n306) );
  NANDX2 U361 ( .IN1(n189), .IN2(n408), .OUT(n303) );
  NANDX2 U362 ( .IN1(n185), .IN2(n380), .OUT(n392) );
  NANDX2 U363 ( .IN1(n356), .IN2(n179), .OUT(n305) );
  INVX4 U364 ( .IN(n358), .OUT(n366) );
  INVX4 U365 ( .IN(n175), .OUT(n227) );
  INVX4 U366 ( .IN(n795), .OUT(n323) );
  NANDX2 U367 ( .IN1(n344), .IN2(n499), .OUT(n795) );
  INVX4 U368 ( .IN(n169), .OUT(n499) );
  NANDX2 U369 ( .IN1(n449), .IN2(n233), .OUT(n448) );
  NANDX2 U370 ( .IN1(n441), .IN2(n226), .OUT(n449) );
  NANDX2 U371 ( .IN1(Multi_dataout[2]), .IN2(n231), .OUT(n441) );
  NANDX2 U372 ( .IN1(n205), .IN2(n482), .OUT(n446) );
  NANDX2 U373 ( .IN1(n217), .IN2(n482), .OUT(n406) );
  INVX4 U374 ( .IN(n204), .OUT(n482) );
  INVX4 U375 ( .IN(n312), .OUT(n407) );
  NANDX2 U376 ( .IN1(n184), .IN2(n386), .OUT(n430) );
  NANDX2 U377 ( .IN1(n183), .IN2(n187), .OUT(n386) );
  INVX4 U378 ( .IN(n429), .OUT(n187) );
  NANDX2 U379 ( .IN1(n178), .IN2(n378), .OUT(n429) );
  NANDX2 U380 ( .IN1(n177), .IN2(n178), .OUT(n378) );
  NANDX2 U381 ( .IN1(n176), .IN2(n509), .OUT(n177) );
  INVX4 U382 ( .IN(Multi_dataout[11]), .OUT(n509) );
  INVX4 U383 ( .IN(n410), .OUT(n178) );
  NANDX2 U384 ( .IN1(n455), .IN2(n508), .OUT(n410) );
  NANDX2 U385 ( .IN1(n182), .IN2(n510), .OUT(n183) );
  INVX4 U386 ( .IN(Multi_dataout[9]), .OUT(n510) );
  INVX4 U387 ( .IN(n167), .OUT(n502) );
  INVX4 U388 ( .IN(n789), .OUT(n344) );
  INVX4 U389 ( .IN(n281), .OUT(n289) );
  INVX4 U390 ( .IN(n278), .OUT(n272) );
  NAND2X1 U391 ( .IN1(RSTn), .IN2(n861), .OUT(n320) );
  INVX4 U392 ( .IN(Multi_ack), .OUT(n836) );
  INVX4 U393 ( .IN(n604), .OUT(Dataout_valid) );
  INVX1 U394 ( .IN(n433), .OUT(n434) );
  INVX1 U395 ( .IN(n783), .OUT(n767) );
  NAND2X1 U396 ( .IN1(n397), .IN2(n402), .OUT(n398) );
  NAND2X1 U397 ( .IN1(n397), .IN2(n400), .OUT(n396) );
  INVX1 U398 ( .IN(n798), .OUT(n862) );
  NAND2X1 U399 ( .IN1(n465), .IN2(n415), .OUT(n416) );
  NAND2X1 U400 ( .IN1(Debug_reg[1]), .IN2(n411), .OUT(n414) );
  BUF4X U401 ( .IN(n758), .OUT(n114) );
  BUF4X U402 ( .IN(n757), .OUT(n113) );
  INVX1 U403 ( .IN(n372), .OUT(n374) );
  INVX1 U404 ( .IN(n545), .OUT(n550) );
  INVX1 U405 ( .IN(n246), .OUT(n247) );
  NAND2X1 U406 ( .IN1(n109), .IN2(n279), .OUT(n242) );
  NAND2X1 U407 ( .IN1(Datain1[9]), .IN2(n497), .OUT(n259) );
  INVX1 U408 ( .IN(n271), .OUT(n287) );
  INVX1 U409 ( .IN(n267), .OUT(n283) );
  INVX1 U410 ( .IN(n330), .OUT(n286) );
  NAND2X1 U411 ( .IN1(Final_Exponent_reg[5]), .IN2(n647), .OUT(n274) );
  NAND2X1 U412 ( .IN1(n278), .IN2(n279), .OUT(n273) );
  INVX1 U413 ( .IN(n111), .OUT(DP_OP_433J3_126_901_n15) );
  NAND2X1 U414 ( .IN1(n337), .IN2(n336), .OUT(n338) );
  INVX1 U415 ( .IN(n501), .OUT(n241) );
  INVX1 U416 ( .IN(n644), .OUT(n331) );
  NAND2X1 U417 ( .IN1(n465), .IN2(n464), .OUT(n466) );
  INVX1 U418 ( .IN(n365), .OUT(n431) );
  NAND2X1 U419 ( .IN1(n455), .IN2(n454), .OUT(n456) );
  INVX1 U420 ( .IN(n352), .OUT(n353) );
  NAND2X1 U421 ( .IN1(n465), .IN2(n408), .OUT(n445) );
  NAND2X1 U422 ( .IN1(n465), .IN2(n427), .OUT(n428) );
  INVX4 U423 ( .IN(n481), .OUT(n465) );
  INVX1 U424 ( .IN(Mode[1]), .OUT(n403) );
  INVX1 U425 ( .IN(Mode[0]), .OUT(n506) );
  NAND2X1 U426 ( .IN1(Datain2[8]), .IN2(n530), .OUT(n83) );
  NAND2X1 U427 ( .IN1(Datain1[8]), .IN2(n524), .OUT(n82) );
  INVX1 U428 ( .IN(n619), .OUT(n143) );
  NAND2X1 U429 ( .IN1(Datain2[9]), .IN2(n529), .OUT(n87) );
  NAND2X1 U430 ( .IN1(Datain1[9]), .IN2(n85), .OUT(n86) );
  INVX1 U431 ( .IN(Datain2[9]), .OUT(n85) );
  NAND2X1 U432 ( .IN1(Datain2[10]), .IN2(n89), .OUT(n91) );
  NAND2X1 U433 ( .IN1(Datain1[10]), .IN2(n520), .OUT(n90) );
  NAND2X1 U434 ( .IN1(Datain2[11]), .IN2(n533), .OUT(n95) );
  NAND2X1 U435 ( .IN1(Datain1[11]), .IN2(n521), .OUT(n93) );
  NAND2X1 U436 ( .IN1(Datain2[12]), .IN2(n532), .OUT(n100) );
  NAND2X1 U437 ( .IN1(Datain1[12]), .IN2(n98), .OUT(n99) );
  INVX1 U438 ( .IN(Datain2[12]), .OUT(n98) );
  NAND2X1 U439 ( .IN1(Datain2[13]), .IN2(n103), .OUT(n105) );
  INVX1 U440 ( .IN(Datain1[13]), .OUT(n103) );
  NAND2X1 U441 ( .IN1(Datain1[13]), .IN2(n102), .OUT(n104) );
  INVX1 U442 ( .IN(Datain2[13]), .OUT(n102) );
  NAND2X1 U443 ( .IN1(n58), .IN2(n227), .OUT(n221) );
  NAND2X1 U444 ( .IN1(n358), .IN2(n209), .OUT(n210) );
  NAND2X1 U445 ( .IN1(n358), .IN2(n367), .OUT(n219) );
  NAND2X1 U446 ( .IN1(Multi_dataout[8]), .IN2(n510), .OUT(n197) );
  NAND2X1 U447 ( .IN1(Multi_dataout[10]), .IN2(n509), .OUT(n191) );
  NAND2X1 U448 ( .IN1(n642), .IN2(n360), .OUT(n192) );
  NAND2X1 U449 ( .IN1(n644), .IN2(n366), .OUT(n189) );
  NAND2X1 U450 ( .IN1(n116), .IN2(Final_Exponent_reg[2]), .OUT(n180) );
  INVX1 U451 ( .IN(Multi_dataout[4]), .OUT(n211) );
  INVX1 U452 ( .IN(Multi_dataout[5]), .OUT(n212) );
  NAND2X1 U453 ( .IN1(Multi_dataout[6]), .IN2(n187), .OUT(n188) );
  INVX1 U454 ( .IN(Multi_dataout[7]), .OUT(n181) );
  INVX1 U455 ( .IN(Multi_dataout[8]), .OUT(n182) );
  BUF4X U456 ( .IN(Final_Exponent_reg[1]), .OUT(n116) );
  INVX1 U457 ( .IN(Datain1[10]), .OUT(n89) );
  TIEHI U458 ( .OUT(n64) );
  NAND2X1 U459 ( .IN1(Multi_dataout[11]), .IN2(n178), .OUT(n454) );
  NAND2X1 U460 ( .IN1(Multi_dataout[12]), .IN2(n455), .OUT(n354) );
  INVX1 U461 ( .IN(n108), .OUT(DP_OP_433J3_126_901_n23) );
  INVX1 U462 ( .IN(C1_Z_0), .OUT(n119) );
  INVX1 U463 ( .IN(n386), .OUT(n409) );
  BUF4X U464 ( .IN(n410), .OUT(n110) );
  INVX1 U465 ( .IN(n406), .OUT(n218) );
  NAND2X1 U466 ( .IN1(n412), .IN2(n446), .OUT(n413) );
  INVX1 U467 ( .IN(n446), .OUT(n382) );
  INVX1 U468 ( .IN(n314), .OUT(n442) );
  NAND2X1 U469 ( .IN1(n465), .IN2(n429), .OUT(n438) );
  INVX1 U470 ( .IN(n412), .OUT(n367) );
  NAND2X1 U471 ( .IN1(n442), .IN2(n441), .OUT(n443) );
  NAND2X1 U472 ( .IN1(n431), .IN2(n430), .OUT(n432) );
  NAND2X1 U473 ( .IN1(n378), .IN2(n430), .OUT(n312) );
  NAND2X1 U474 ( .IN1(n386), .IN2(n430), .OUT(n437) );
  INVX1 U475 ( .IN(n231), .OUT(n224) );
  INVX1 U476 ( .IN(Multi_dataout[12]), .OUT(n508) );
  INVX1 U477 ( .IN(DP_OP_433J3_126_901_n11), .OUT(n121) );
  INVX1 U478 ( .IN(DP_OP_433J3_126_901_n7), .OUT(n122) );
  INVX4 U479 ( .IN(n635), .OUT(n583) );
  INVX4 U480 ( .IN(n779), .OUT(n579) );
  NOR2X1 U481 ( .IN1(n526), .IN2(n525), .OUT(n619) );
  NOR2X1 U482 ( .IN1(n535), .IN2(n534), .OUT(n618) );
  INVX4 U483 ( .IN(n777), .OUT(n504) );
  NOR2X1 U484 ( .IN1(n53), .IN2(n709), .OUT(n164) );
  AOI21 U485 ( .IN1(N392), .IN2(n504), .IN3(n165), .OUT(n545) );
  INVX4 U486 ( .IN(n585), .OUT(n503) );
  NANDX2 U487 ( .IN1(n503), .IN2(Multi_ack), .OUT(n794) );
  MUX2X1 U488 ( .IN1(n60), .IN2(Final_Exponent_reg[8]), .S(n288), .OUT(n492)
         );
  INVX4 U489 ( .IN(n632), .OUT(n511) );
  NOR2X1 U490 ( .IN1(n772), .IN2(StateMC[0]), .OUT(n778) );
  AOI21 U491 ( .IN1(n503), .IN2(n640), .IN3(n861), .OUT(n330) );
  OAI21 U492 ( .IN1(n126), .IN2(n330), .IN3(n884), .OUT(n293) );
  INVX4 U493 ( .IN(n385), .OUT(n486) );
  NOR2X1 U494 ( .IN1(Final_Exponent_reg[4]), .IN2(Final_Exponent_reg[6]), 
        .OUT(n174) );
  NOR2X1 U495 ( .IN1(Final_Exponent_reg[7]), .IN2(Final_Exponent_reg[5]), 
        .OUT(n173) );
  NAND3X1 U496 ( .IN1(n60), .IN2(n174), .IN3(n173), .OUT(n175) );
  NOR2X1 U497 ( .IN1(n510), .IN2(n429), .OUT(n365) );
  NOR2X1 U498 ( .IN1(n181), .IN2(n429), .OUT(n184) );
  NAND3X1 U499 ( .IN1(n393), .IN2(n305), .IN3(n392), .OUT(n208) );
  NOR2X1 U500 ( .IN1(n188), .IN2(n437), .OUT(n408) );
  OAI21 U501 ( .IN1(Final_Exponent_reg[0]), .IN2(n356), .IN3(n190), .OUT(n193)
         );
  NOR2X1 U502 ( .IN1(n191), .IN2(n110), .OUT(n352) );
  NOR2X1 U503 ( .IN1(n197), .IN2(n429), .OUT(n427) );
  NOR2X1 U504 ( .IN1(n116), .IN2(Final_Exponent_reg[2]), .OUT(n199) );
  OAI21 U505 ( .IN1(Final_Exponent_reg[0]), .IN2(n209), .IN3(n358), .OUT(n381)
         );
  NOR2X1 U506 ( .IN1(Multi_dataout[6]), .IN2(n429), .OUT(n201) );
  NOR2X1 U507 ( .IN1(n381), .IN2(n446), .OUT(n294) );
  NOR2X1 U508 ( .IN1(n206), .IN2(n294), .OUT(n207) );
  NOR2X1 U509 ( .IN1(n208), .IN2(n372), .OUT(n236) );
  NAND3X1 U510 ( .IN1(Multi_dataout[3]), .IN2(n212), .IN3(n211), .OUT(n216) );
  OAI21 U511 ( .IN1(n642), .IN2(n59), .IN3(n390), .OUT(n223) );
  NOR2X1 U512 ( .IN1(n222), .IN2(n314), .OUT(n231) );
  NOR2X1 U513 ( .IN1(n225), .IN2(n224), .OUT(n226) );
  NAND3X1 U514 ( .IN1(n231), .IN2(Multi_dataout[0]), .IN3(n441), .OUT(n232) );
  NOR2X1 U515 ( .IN1(n235), .IN2(n300), .OUT(n495) );
  INVX4 U516 ( .IN(n237), .OUT(n339) );
  AOI22 U517 ( .IN1(n498), .IN2(Datain2[7]), .IN3(n497), .IN4(Datain1[7]), 
        .OUT(n244) );
  INVX4 U518 ( .IN(n596), .OUT(n500) );
  NOR2X1 U519 ( .IN1(n512), .IN2(n639), .OUT(n501) );
  NAND3X1 U520 ( .IN1(n244), .IN2(n243), .IN3(n242), .OUT(n245) );
  AOI21 U521 ( .IN1(C276_DATA3_0), .IN2(n339), .IN3(n245), .OUT(n246) );
  AOI22 U522 ( .IN1(Final_Exponent_reg[0]), .IN2(n293), .IN3(RSTn), .IN4(n247), 
        .OUT(n250) );
  NOR2X1 U523 ( .IN1(n628), .IN2(n660), .OUT(n267) );
  AOI22 U524 ( .IN1(n492), .IN2(n501), .IN3(n500), .IN4(N392), .OUT(n345) );
  INVX4 U525 ( .IN(n340), .OUT(n266) );
  AOI21 U526 ( .IN1(n109), .IN2(n116), .IN3(n641), .OUT(n252) );
  AOI22 U527 ( .IN1(n498), .IN2(Datain2[8]), .IN3(n497), .IN4(Datain1[8]), 
        .OUT(n251) );
  OAI21 U528 ( .IN1(n252), .IN2(n649), .IN3(n251), .OUT(n253) );
  AOI21 U529 ( .IN1(n500), .IN2(N385), .IN3(n253), .OUT(n255) );
  AOI22 U530 ( .IN1(n116), .IN2(n293), .IN3(RSTn), .IN4(n256), .OUT(n257) );
  AOI22 U531 ( .IN1(n643), .IN2(n58), .IN3(Datain2[9]), .IN4(n498), .OUT(n260)
         );
  NAND3X1 U532 ( .IN1(n55), .IN2(n642), .IN3(n279), .OUT(n258) );
  NAND3X1 U533 ( .IN1(n260), .IN2(n259), .IN3(n258), .OUT(n261) );
  AOI21 U534 ( .IN1(N386), .IN2(n500), .IN3(n261), .OUT(n263) );
  AOI22 U535 ( .IN1(n55), .IN2(n293), .IN3(RSTn), .IN4(n264), .OUT(n265) );
  AOI22 U536 ( .IN1(n498), .IN2(Datain2[11]), .IN3(n497), .IN4(Datain1[11]), 
        .OUT(n270) );
  AOI22 U537 ( .IN1(n648), .IN2(n71), .IN3(n330), .IN4(n273), .OUT(n268) );
  AOI22 U538 ( .IN1(n498), .IN2(Datain2[12]), .IN3(n497), .IN4(Datain1[12]), 
        .OUT(n276) );
  NAND3X1 U539 ( .IN1(n272), .IN2(n69), .IN3(n279), .OUT(n275) );
  NAND3X1 U540 ( .IN1(n276), .IN2(n275), .IN3(n274), .OUT(n277) );
  AOI22 U541 ( .IN1(n498), .IN2(Datain2[13]), .IN3(n497), .IN4(Datain1[13]), 
        .OUT(n284) );
  OAI21 U542 ( .IN1(n69), .IN2(n278), .IN3(n75), .OUT(n280) );
  NAND3X1 U543 ( .IN1(n281), .IN2(n280), .IN3(n279), .OUT(n282) );
  NAND3X1 U544 ( .IN1(n284), .IN2(n283), .IN3(n282), .OUT(n285) );
  OAI21 U545 ( .IN1(Final_Exponent_reg[7]), .IN2(n289), .IN3(n288), .OUT(n291)
         );
  AOI22 U546 ( .IN1(n498), .IN2(Datain2[14]), .IN3(n497), .IN4(Datain1[14]), 
        .OUT(n290) );
  OAI21 U547 ( .IN1(n291), .IN2(n649), .IN3(n290), .OUT(n292) );
  NAND3X1 U548 ( .IN1(n298), .IN2(n394), .IN3(n310), .OUT(C1_Z_3) );
  NAND3X1 U549 ( .IN1(n392), .IN2(n393), .IN3(n650), .OUT(n301) );
  NOR2X1 U550 ( .IN1(n301), .IN2(n300), .OUT(n302) );
  NAND3X1 U551 ( .IN1(n306), .IN2(n305), .IN3(n304), .OUT(n307) );
  NOR2X1 U552 ( .IN1(n308), .IN2(n307), .OUT(n309) );
  NAND3X1 U553 ( .IN1(n311), .IN2(n650), .IN3(n310), .OUT(C1_Z_0) );
  NAND3X1 U554 ( .IN1(n386), .IN2(n354), .IN3(n407), .OUT(n313) );
  NOR2X1 U555 ( .IN1(n313), .IN2(n408), .OUT(n315) );
  NOR2X1 U556 ( .IN1(n460), .IN2(n464), .OUT(n433) );
  NAND3X1 U557 ( .IN1(n452), .IN2(n884), .IN3(n320), .OUT(n328) );
  AOI22 U558 ( .IN1(n492), .IN2(n502), .IN3(Final_Exponent_reg[8]), .IN4(n321), 
        .OUT(n325) );
  NAND3X1 U559 ( .IN1(n323), .IN2(n322), .IN3(C276_DATA3_8), .OUT(n324) );
  OAI21 U560 ( .IN1(n794), .IN2(n326), .IN3(n345), .OUT(n327) );
  AOI22 U561 ( .IN1(Final_Exponent_reg[8]), .IN2(n328), .IN3(RSTn), .IN4(n327), 
        .OUT(n329) );
  OAI21 U562 ( .IN1(n331), .IN2(n649), .IN3(n330), .OUT(n335) );
  AOI22 U563 ( .IN1(n645), .IN2(n59), .IN3(Datain2[10]), .IN4(n498), .OUT(n332) );
  OAI21 U564 ( .IN1(n333), .IN2(n89), .IN3(n332), .OUT(n334) );
  AOI21 U565 ( .IN1(n335), .IN2(Final_Exponent_reg[3]), .IN3(n334), .OUT(n337)
         );
  AOI21 U566 ( .IN1(C276_DATA3_3), .IN2(n339), .IN3(n338), .OUT(n342) );
  AOI21 U567 ( .IN1(Final_Exponent_reg[3]), .IN2(n496), .IN3(n340), .OUT(n341)
         );
  OAI21 U568 ( .IN1(n126), .IN2(n342), .IN3(n341), .OUT(n876) );
  NAND3X1 U569 ( .IN1(Mode[2]), .IN2(Mode[1]), .IN3(n506), .OUT(n420) );
  OAI21 U570 ( .IN1(n596), .IN2(N392), .IN3(n609), .OUT(n343) );
  AOI22 U571 ( .IN1(n598), .IN2(Exc_value[2]), .IN3(n74), .IN4(n343), .OUT(
        n591) );
  NAND3X1 U572 ( .IN1(n602), .IN2(n603), .IN3(n345), .OUT(n606) );
  OAI21 U573 ( .IN1(n777), .IN2(N392), .IN3(n609), .OUT(n348) );
  AOI21 U574 ( .IN1(n348), .IN2(n80), .IN3(n347), .OUT(n617) );
  NANDX2 U575 ( .IN1(RSTn), .IN2(n504), .OUT(n349) );
  OAI21 U576 ( .IN1(n59), .IN2(n433), .IN3(n350), .OUT(n351) );
  OAI21 U577 ( .IN1(n356), .IN2(n454), .IN3(n355), .OUT(n357) );
  NOR2X1 U578 ( .IN1(n357), .IN2(n427), .OUT(n362) );
  NOR2X1 U579 ( .IN1(n116), .IN2(n358), .OUT(n359) );
  OAI21 U580 ( .IN1(n360), .IN2(n359), .IN3(n380), .OUT(n361) );
  NOR2X1 U581 ( .IN1(n363), .IN2(n406), .OUT(n387) );
  NOR2X1 U582 ( .IN1(n364), .IN2(n387), .OUT(n370) );
  AOI21 U583 ( .IN1(n367), .IN2(n366), .IN3(n408), .OUT(n389) );
  OAI21 U584 ( .IN1(n368), .IN2(n431), .IN3(n389), .OUT(n369) );
  AOI21 U585 ( .IN1(n415), .IN2(n390), .IN3(n369), .OUT(n384) );
  OAI21 U586 ( .IN1(n464), .IN2(n371), .IN3(Final_Exponent_reg[0]), .OUT(n377)
         );
  NAND3X1 U587 ( .IN1(n374), .IN2(n373), .IN3(n395), .OUT(n375) );
  AOI21 U588 ( .IN1(n382), .IN2(n381), .IN3(n380), .OUT(n388) );
  NOR2X1 U589 ( .IN1(n782), .IN2(n385), .OUT(n397) );
  AOI21 U590 ( .IN1(n754), .IN2(n755), .IN3(n753), .OUT(n401) );
  MUX2X1 U591 ( .IN1(n401), .IN2(n756), .S(n400), .OUT(n783) );
  MUX2X1 U592 ( .IN1(n787), .IN2(n788), .S(n402), .OUT(n791) );
  AOI21 U593 ( .IN1(n491), .IN2(n420), .IN3(n832), .OUT(n489) );
  NOR2X1 U594 ( .IN1(n855), .IN2(n857), .OUT(n426) );
  AOI21 U595 ( .IN1(n405), .IN2(n465), .IN3(n404), .OUT(n424) );
  NAND3X1 U596 ( .IN1(n407), .IN2(n406), .IN3(n441), .OUT(n418) );
  OAI21 U597 ( .IN1(n110), .IN2(n409), .IN3(n465), .OUT(n411) );
  AOI22 U598 ( .IN1(n445), .IN2(n414), .IN3(n465), .IN4(n413), .OUT(n417) );
  AOI22 U599 ( .IN1(n465), .IN2(n418), .IN3(n417), .IN4(n416), .OUT(n419) );
  AOI22 U600 ( .IN1(n424), .IN2(n423), .IN3(n422), .IN4(N392), .OUT(n425) );
  OAI21 U601 ( .IN1(n483), .IN2(n426), .IN3(n425), .OUT(n797) );
  NAND3X1 U602 ( .IN1(Debug_reg[3]), .IN2(n438), .IN3(n457), .OUT(n435) );
  OAI21 U603 ( .IN1(n453), .IN2(n435), .IN3(n480), .OUT(n436) );
  AOI21 U604 ( .IN1(Debug_reg[2]), .IN2(n438), .IN3(n437), .OUT(n439) );
  OAI21 U605 ( .IN1(n465), .IN2(Debug_reg[2]), .IN3(n440), .OUT(n444) );
  AOI22 U606 ( .IN1(n445), .IN2(n444), .IN3(n465), .IN4(n443), .OUT(n451) );
  OAI21 U607 ( .IN1(n481), .IN2(n446), .IN3(n451), .OUT(n447) );
  NAND3X1 U608 ( .IN1(n449), .IN2(n448), .IN3(n447), .OUT(n450) );
  OAI21 U609 ( .IN1(n465), .IN2(n451), .IN3(n450), .OUT(n827) );
  OAI21 U610 ( .IN1(n69), .IN2(n581), .IN3(n568), .OUT(ExcCheck_Datain[12]) );
  OAI21 U611 ( .IN1(n75), .IN2(n581), .IN3(n569), .OUT(ExcCheck_Datain[13]) );
  OAI21 U612 ( .IN1(n72), .IN2(n581), .IN3(n570), .OUT(ExcCheck_Datain[14]) );
  AOI21 U613 ( .IN1(n456), .IN2(n465), .IN3(n468), .OUT(n458) );
  AOI22 U614 ( .IN1(n465), .IN2(n459), .IN3(n458), .IN4(n457), .OUT(n461) );
  AOI22 U615 ( .IN1(n462), .IN2(n461), .IN3(n465), .IN4(n460), .OUT(n463) );
  NOR2X1 U616 ( .IN1(n795), .IN2(n463), .OUT(n467) );
  AOI22 U617 ( .IN1(n795), .IN2(n468), .IN3(n467), .IN4(n466), .OUT(n470) );
  OAI21 U618 ( .IN1(n490), .IN2(n470), .IN3(n469), .OUT(n471) );
  OAI21 U619 ( .IN1(n474), .IN2(n473), .IN3(n472), .OUT(n475) );
  OAI21 U620 ( .IN1(RSOP_428_C1_Z_0), .IN2(n484), .IN3(n475), .OUT(n476) );
  AOI22 U621 ( .IN1(Debug_reg[0]), .IN2(n477), .IN3(RSTn), .IN4(n476), .OUT(
        n478) );
  AOI22 U622 ( .IN1(Debug_reg[0]), .IN2(n563), .IN3(StateMC[0]), .IN4(n562), 
        .OUT(n479) );
  NOR2X1 U623 ( .IN1(n69), .IN2(n604), .OUT(Dataout[12]) );
  NOR2X1 U624 ( .IN1(n75), .IN2(n604), .OUT(Dataout[13]) );
  NOR2X1 U625 ( .IN1(n72), .IN2(n604), .OUT(Dataout[14]) );
  OAI21 U626 ( .IN1(n482), .IN2(n481), .IN3(n480), .OUT(n487) );
  AOI21 U627 ( .IN1(n487), .IN2(n486), .IN3(n485), .OUT(n488) );
  NOR2X1 U628 ( .IN1(n126), .IN2(n488), .OUT(n96) );
  NAND3X1 U629 ( .IN1(StateMC[2]), .IN2(n66), .IN3(n57), .OUT(n635) );
  NOR2X1 U630 ( .IN1(n214), .IN2(n215), .OUT(n513) );
  NAND3X1 U631 ( .IN1(Exc_value[0]), .IN2(Exc_value[1]), .IN3(n513), .OUT(n601) );
  INVX1 U632 ( .IN(Exc_value[2]), .OUT(n599) );
  NOR2X1 U633 ( .IN1(n599), .IN2(n213), .OUT(n515) );
  INVX1 U634 ( .IN(Exc_value[0]), .OUT(n613) );
  NAND2X1 U635 ( .IN1(Exc_value[2]), .IN2(n613), .OUT(n514) );
  NOR2X1 U636 ( .IN1(Exc_value[1]), .IN2(n514), .OUT(n634) );
  OAI21 U637 ( .IN1(n601), .IN2(n515), .IN3(n630), .OUT(n636) );
  NAND2X1 U638 ( .IN1(StateMC[2]), .IN2(n57), .OUT(n516) );
  NOR2X1 U639 ( .IN1(n66), .IN2(n516), .OUT(n709) );
  NAND3X1 U640 ( .IN1(Datain1[10]), .IN2(Datain1[13]), .IN3(Datain1[11]), 
        .OUT(n517) );
  NOR2X1 U641 ( .IN1(n529), .IN2(n517), .OUT(n518) );
  NAND3X1 U642 ( .IN1(Datain1[7]), .IN2(Datain1[12]), .IN3(n518), .OUT(n527)
         );
  NOR2X1 U643 ( .IN1(Datain2[9]), .IN2(Datain2[13]), .OUT(n519) );
  NAND3X1 U644 ( .IN1(n521), .IN2(n520), .IN3(n519), .OUT(n526) );
  NOR2X1 U645 ( .IN1(Datain2[14]), .IN2(Datain2[12]), .OUT(n522) );
  NAND3X1 U646 ( .IN1(n524), .IN2(n523), .IN3(n522), .OUT(n525) );
  OAI21 U647 ( .IN1(n530), .IN2(n527), .IN3(n619), .OUT(n542) );
  NOR2X1 U648 ( .IN1(Datain1[13]), .IN2(Datain1[10]), .OUT(n528) );
  NAND3X1 U649 ( .IN1(n530), .IN2(n529), .IN3(n528), .OUT(n535) );
  NOR2X1 U650 ( .IN1(Datain1[14]), .IN2(Datain1[7]), .OUT(n531) );
  NAND3X1 U651 ( .IN1(n533), .IN2(n532), .IN3(n531), .OUT(n534) );
  INVX1 U652 ( .IN(Datain2[14]), .OUT(n540) );
  NAND2X1 U653 ( .IN1(Datain2[10]), .IN2(Datain2[11]), .OUT(n537) );
  NAND3X1 U654 ( .IN1(Datain2[13]), .IN2(Datain2[8]), .IN3(Datain2[9]), .OUT(
        n536) );
  NOR2X1 U655 ( .IN1(n537), .IN2(n536), .OUT(n538) );
  NAND3X1 U656 ( .IN1(Datain2[12]), .IN2(Datain2[7]), .IN3(n538), .OUT(n539)
         );
  NAND3X1 U657 ( .IN1(n618), .IN2(n540), .IN3(n539), .OUT(n541) );
  OAI21 U658 ( .IN1(Datain1[14]), .IN2(n542), .IN3(n541), .OUT(n610) );
  NAND3X1 U659 ( .IN1(n545), .IN2(n794), .IN3(n544), .OUT(n546) );
  AOI21 U660 ( .IN1(n583), .IN2(n636), .IN3(n546), .OUT(n547) );
  NAND3X1 U661 ( .IN1(StateMC[1]), .IN2(StateMC[0]), .IN3(n65), .OUT(n779) );
  AOI21 U662 ( .IN1(n547), .IN2(n629), .IN3(n126), .OUT(N90) );
  NOR2X1 U663 ( .IN1(n59), .IN2(n644), .OUT(n646) );
  AOI21 U664 ( .IN1(Multi_dataout[15]), .IN2(n492), .IN3(n789), .OUT(n549) );
  AOI22 U665 ( .IN1(n579), .IN2(n548), .IN3(n778), .IN4(Data_valid), .OUT(n553) );
  OAI21 U666 ( .IN1(n549), .IN2(n794), .IN3(n553), .OUT(n551) );
  NOR2X1 U667 ( .IN1(n551), .IN2(n550), .OUT(n552) );
  AOI21 U668 ( .IN1(n552), .IN2(n632), .IN3(n126), .OUT(N89) );
  AOI21 U669 ( .IN1(n52), .IN2(n53), .IN3(n504), .OUT(n555) );
  NAND2X1 U670 ( .IN1(G_reg), .IN2(Final_Mantissa_reg[0]), .OUT(n674) );
  NOR2X1 U671 ( .IN1(n674), .IN2(n62), .OUT(n693) );
  NOR2X1 U672 ( .IN1(n63), .IN2(n707), .OUT(n728) );
  NOR2X1 U673 ( .IN1(n740), .IN2(n67), .OUT(n748) );
  AOI22 U674 ( .IN1(n501), .IN2(n492), .IN3(n511), .IN4(n636), .OUT(n554) );
  NAND3X1 U675 ( .IN1(n555), .IN2(n554), .IN3(n585), .OUT(n556) );
  OAI21 U676 ( .IN1(n557), .IN2(n556), .IN3(RSTn), .OUT(n703) );
  NOR2X1 U677 ( .IN1(n76), .IN2(n604), .OUT(Dataout[0]) );
  NOR2X1 U678 ( .IN1(n59), .IN2(n604), .OUT(Dataout[10]) );
  NOR2X1 U679 ( .IN1(n71), .IN2(n604), .OUT(Dataout[11]) );
  NOR2X1 U680 ( .IN1(n604), .IN2(n78), .OUT(Dataout[15]) );
  NOR2X1 U681 ( .IN1(n62), .IN2(n604), .OUT(Dataout[1]) );
  NOR2X1 U682 ( .IN1(n70), .IN2(n604), .OUT(Dataout[2]) );
  NOR2X1 U683 ( .IN1(n63), .IN2(n604), .OUT(Dataout[3]) );
  NOR2X1 U684 ( .IN1(n68), .IN2(n604), .OUT(Dataout[4]) );
  NOR2X1 U685 ( .IN1(n67), .IN2(n604), .OUT(Dataout[5]) );
  NOR2X1 U686 ( .IN1(n73), .IN2(n604), .OUT(Dataout[6]) );
  NOR2X1 U687 ( .IN1(n109), .IN2(n604), .OUT(Dataout[7]) );
  NOR2X1 U688 ( .IN1(n61), .IN2(n604), .OUT(Dataout[8]) );
  NOR2X1 U689 ( .IN1(n58), .IN2(n604), .OUT(Dataout[9]) );
  NAND2X1 U690 ( .IN1(Mode[2]), .IN2(n506), .OUT(n558) );
  NOR2X1 U691 ( .IN1(Mode[1]), .IN2(n558), .OUT(n562) );
  AOI22 U692 ( .IN1(StateMC[1]), .IN2(n562), .IN3(Debug_reg[1]), .IN4(n563), 
        .OUT(n559) );
  AOI22 U693 ( .IN1(StateMC[2]), .IN2(n562), .IN3(Debug_reg[2]), .IN4(n563), 
        .OUT(n560) );
  NAND2X1 U694 ( .IN1(n563), .IN2(Debug_reg[3]), .OUT(n561) );
  AOI21 U695 ( .IN1(Debug_valid_reg), .IN2(n563), .IN3(n562), .OUT(n564) );
  AOI22 U696 ( .IN1(n579), .IN2(Datain1[0]), .IN3(n583), .IN4(Datain2[0]), 
        .OUT(n565) );
  OAI21 U697 ( .IN1(n76), .IN2(n581), .IN3(n565), .OUT(ExcCheck_Datain[0]) );
  AOI22 U698 ( .IN1(n579), .IN2(Datain1[10]), .IN3(Datain2[10]), .IN4(n583), 
        .OUT(n566) );
  OAI21 U699 ( .IN1(n59), .IN2(n581), .IN3(n566), .OUT(ExcCheck_Datain[10]) );
  AOI22 U700 ( .IN1(n579), .IN2(Datain1[11]), .IN3(Datain2[11]), .IN4(n583), 
        .OUT(n567) );
  OAI21 U701 ( .IN1(n71), .IN2(n581), .IN3(n567), .OUT(ExcCheck_Datain[11]) );
  AOI22 U702 ( .IN1(n579), .IN2(Datain1[12]), .IN3(Datain2[12]), .IN4(n583), 
        .OUT(n568) );
  AOI22 U703 ( .IN1(n579), .IN2(Datain1[13]), .IN3(Datain2[13]), .IN4(n583), 
        .OUT(n569) );
  AOI22 U704 ( .IN1(n579), .IN2(Datain1[14]), .IN3(Datain2[14]), .IN4(n583), 
        .OUT(n570) );
  AOI22 U705 ( .IN1(n579), .IN2(Datain1[1]), .IN3(n583), .IN4(Datain2[1]), 
        .OUT(n571) );
  OAI21 U706 ( .IN1(n62), .IN2(n581), .IN3(n571), .OUT(ExcCheck_Datain[1]) );
  AOI22 U707 ( .IN1(n579), .IN2(Datain1[2]), .IN3(n583), .IN4(Datain2[2]), 
        .OUT(n572) );
  OAI21 U708 ( .IN1(n70), .IN2(n581), .IN3(n572), .OUT(ExcCheck_Datain[2]) );
  AOI22 U709 ( .IN1(n579), .IN2(Datain1[3]), .IN3(n583), .IN4(Datain2[3]), 
        .OUT(n573) );
  OAI21 U710 ( .IN1(n63), .IN2(n581), .IN3(n573), .OUT(ExcCheck_Datain[3]) );
  AOI22 U711 ( .IN1(n579), .IN2(Datain1[4]), .IN3(n583), .IN4(Datain2[4]), 
        .OUT(n574) );
  OAI21 U712 ( .IN1(n68), .IN2(n581), .IN3(n574), .OUT(ExcCheck_Datain[4]) );
  AOI22 U713 ( .IN1(n579), .IN2(Datain1[5]), .IN3(n583), .IN4(Datain2[5]), 
        .OUT(n575) );
  OAI21 U714 ( .IN1(n67), .IN2(n581), .IN3(n575), .OUT(ExcCheck_Datain[5]) );
  AOI22 U715 ( .IN1(n579), .IN2(Datain1[6]), .IN3(n583), .IN4(Datain2[6]), 
        .OUT(n576) );
  OAI21 U716 ( .IN1(n73), .IN2(n581), .IN3(n576), .OUT(ExcCheck_Datain[6]) );
  AOI22 U717 ( .IN1(n579), .IN2(Datain1[7]), .IN3(Datain2[7]), .IN4(n583), 
        .OUT(n577) );
  OAI21 U718 ( .IN1(n109), .IN2(n581), .IN3(n577), .OUT(ExcCheck_Datain[7]) );
  AOI22 U719 ( .IN1(n579), .IN2(Datain1[8]), .IN3(Datain2[8]), .IN4(n583), 
        .OUT(n578) );
  OAI21 U720 ( .IN1(n61), .IN2(n581), .IN3(n578), .OUT(ExcCheck_Datain[8]) );
  AOI22 U721 ( .IN1(n579), .IN2(Datain1[9]), .IN3(Datain2[9]), .IN4(n583), 
        .OUT(n580) );
  OAI21 U722 ( .IN1(n58), .IN2(n581), .IN3(n580), .OUT(ExcCheck_Datain[9]) );
  NOR2X1 U723 ( .IN1(n215), .IN2(n604), .OUT(Exc[0]) );
  NOR2X1 U724 ( .IN1(n214), .IN2(n604), .OUT(Exc[1]) );
  NOR2X1 U725 ( .IN1(n213), .IN2(n604), .OUT(Exc[2]) );
  NOR2X1 U726 ( .IN1(T_reg), .IN2(G_reg), .OUT(n594) );
  OAI21 U727 ( .IN1(n628), .IN2(n639), .IN3(n709), .OUT(n582) );
  NOR2X1 U728 ( .IN1(n594), .IN2(n582), .OUT(n615) );
  AOI22 U729 ( .IN1(n634), .IN2(n511), .IN3(n52), .IN4(n584), .OUT(n612) );
  NOR2X1 U730 ( .IN1(n584), .IN2(n583), .OUT(n586) );
  OAI21 U731 ( .IN1(n52), .IN2(n586), .IN3(n585), .OUT(n593) );
  NOR2X1 U732 ( .IN1(n587), .IN2(n593), .OUT(n609) );
  AOI22 U733 ( .IN1(n213), .IN2(Exc_value[2]), .IN3(n599), .IN4(n74), .OUT(
        n588) );
  NOR2X1 U734 ( .IN1(n601), .IN2(n588), .OUT(n589) );
  NAND3X1 U735 ( .IN1(n591), .IN2(n655), .IN3(n590), .OUT(n592) );
  OAI21 U736 ( .IN1(n615), .IN2(n592), .IN3(RSTn), .OUT(n667) );
  NAND3X1 U737 ( .IN1(Multi_dataout[15]), .IN2(n821), .IN3(n492), .OUT(n608)
         );
  AOI21 U738 ( .IN1(n594), .IN2(n709), .IN3(n593), .OUT(n595) );
  AOI22 U739 ( .IN1(Exc_value[1]), .IN2(n598), .IN3(n77), .IN4(n597), .OUT(
        n603) );
  NAND2X1 U740 ( .IN1(n213), .IN2(n599), .OUT(n600) );
  NOR2X1 U741 ( .IN1(n601), .IN2(n600), .OUT(n631) );
  NOR2X1 U742 ( .IN1(n126), .IN2(n604), .OUT(n605) );
  AOI22 U743 ( .IN1(RSTn), .IN2(n606), .IN3(n605), .IN4(n77), .OUT(n607) );
  OAI21 U744 ( .IN1(n854), .IN2(n608), .IN3(n607), .OUT(n883) );
  AOI21 U745 ( .IN1(n511), .IN2(n631), .IN3(Exc[0]), .OUT(n611) );
  OAI21 U746 ( .IN1(n613), .IN2(n612), .IN3(n611), .OUT(n614) );
  NOR2X1 U747 ( .IN1(n615), .IN2(n614), .OUT(n616) );
  AOI21 U748 ( .IN1(n617), .IN2(n616), .IN3(n126), .OUT(n882) );
  NOR2X1 U749 ( .IN1(n126), .IN2(n504), .OUT(n819) );
  AOI21 U750 ( .IN1(n127), .IN2(n619), .IN3(n349), .OUT(n620) );
  AOI21 U751 ( .IN1(Op2_Mantissa_reg[7]), .IN2(n112), .IN3(n620), .OUT(n621)
         );
  OAI21 U752 ( .IN1(Datain2[15]), .IN2(Datain1[15]), .IN3(Data_valid), .OUT(
        n622) );
  AOI21 U753 ( .IN1(Datain2[15]), .IN2(Datain1[15]), .IN3(n622), .OUT(n623) );
  NAND2X1 U754 ( .IN1(RSTn), .IN2(n623), .OUT(n626) );
  NOR2X1 U755 ( .IN1(Data_valid), .IN2(n126), .OUT(n624) );
  OAI21 U756 ( .IN1(n624), .IN2(n627), .IN3(Final_Sign_reg), .OUT(n625) );
  OAI21 U757 ( .IN1(n627), .IN2(n626), .IN3(n625), .OUT(n880) );
  NOR2X1 U758 ( .IN1(n634), .IN2(n631), .OUT(n633) );
  AOI21 U759 ( .IN1(n634), .IN2(n52), .IN3(n779), .OUT(n638) );
  AOI21 U760 ( .IN1(n52), .IN2(n636), .IN3(n635), .OUT(n637) );
  NOR2X1 U761 ( .IN1(n638), .IN2(n637), .OUT(n669) );
  NOR2X1 U762 ( .IN1(n116), .IN2(n109), .OUT(n641) );
  NOR2X1 U763 ( .IN1(n649), .IN2(n642), .OUT(n643) );
  NOR2X1 U764 ( .IN1(n649), .IN2(n644), .OUT(n645) );
  NOR2X1 U765 ( .IN1(n493), .IN2(n494), .OUT(n650) );
  NOR2X1 U766 ( .IN1(n752), .IN2(n754), .OUT(n757) );
  AOI22 U767 ( .IN1(Multi_dataout[2]), .IN2(n716), .IN3(Multi_dataout[1]), 
        .IN4(n113), .OUT(n654) );
  NOR2X1 U768 ( .IN1(n652), .IN2(n752), .OUT(n758) );
  AOI22 U769 ( .IN1(Multi_dataout[3]), .IN2(n717), .IN3(Multi_dataout[0]), 
        .IN4(n114), .OUT(n653) );
  AOI21 U770 ( .IN1(G_reg), .IN2(T_reg), .IN3(Final_Mantissa_reg[0]), .OUT(
        n657) );
  NAND2X1 U771 ( .IN1(n674), .IN2(n709), .OUT(n656) );
  OAI21 U772 ( .IN1(n657), .IN2(n656), .IN3(n655), .OUT(n658) );
  AOI21 U773 ( .IN1(n498), .IN2(Datain2[0]), .IN3(n658), .OUT(n665) );
  NOR2X1 U774 ( .IN1(n781), .IN2(n659), .OUT(n714) );
  AOI22 U775 ( .IN1(Multi_dataout[7]), .IN2(n714), .IN3(n497), .IN4(Datain1[0]), .OUT(n664) );
  NOR2X1 U776 ( .IN1(n492), .IN2(n660), .OUT(n745) );
  AOI22 U777 ( .IN1(Multi_dataout[6]), .IN2(n716), .IN3(Multi_dataout[5]), 
        .IN4(n113), .OUT(n662) );
  AOI22 U778 ( .IN1(Multi_dataout[7]), .IN2(n717), .IN3(Multi_dataout[4]), 
        .IN4(n114), .OUT(n661) );
  AOI22 U779 ( .IN1(Multi_dataout[8]), .IN2(n745), .IN3(n764), .IN4(n733), 
        .OUT(n663) );
  NAND3X1 U780 ( .IN1(n665), .IN2(n664), .IN3(n663), .OUT(n666) );
  AOI21 U781 ( .IN1(n762), .IN2(n725), .IN3(n666), .OUT(n673) );
  AOI21 U782 ( .IN1(n503), .IN2(n668), .IN3(n500), .OUT(n670) );
  AOI21 U783 ( .IN1(n670), .IN2(n669), .IN3(n126), .OUT(n671) );
  NOR2X1 U784 ( .IN1(n496), .IN2(n671), .OUT(n771) );
  NAND2X1 U785 ( .IN1(Final_Mantissa_reg[0]), .IN2(n704), .OUT(n672) );
  OAI21 U786 ( .IN1(n673), .IN2(n126), .IN3(n672), .OUT(n871) );
  AOI21 U787 ( .IN1(n674), .IN2(n62), .IN3(n693), .OUT(n675) );
  AOI22 U788 ( .IN1(Multi_dataout[8]), .IN2(n714), .IN3(n709), .IN4(n675), 
        .OUT(n677) );
  AOI22 U789 ( .IN1(Multi_dataout[9]), .IN2(n745), .IN3(n498), .IN4(Datain2[1]), .OUT(n676) );
  AOI21 U790 ( .IN1(Datain1[1]), .IN2(n497), .IN3(n678), .OUT(n686) );
  AOI22 U791 ( .IN1(Multi_dataout[7]), .IN2(n716), .IN3(Multi_dataout[6]), 
        .IN4(n113), .OUT(n680) );
  AOI22 U792 ( .IN1(Multi_dataout[8]), .IN2(n717), .IN3(Multi_dataout[5]), 
        .IN4(n114), .OUT(n679) );
  AOI22 U793 ( .IN1(Multi_dataout[3]), .IN2(n716), .IN3(Multi_dataout[2]), 
        .IN4(n113), .OUT(n682) );
  AOI22 U794 ( .IN1(Multi_dataout[4]), .IN2(n717), .IN3(Multi_dataout[1]), 
        .IN4(n114), .OUT(n681) );
  AOI22 U795 ( .IN1(n764), .IN2(n743), .IN3(n762), .IN4(n742), .OUT(n685) );
  NOR2X1 U796 ( .IN1(n755), .IN2(n683), .OUT(n741) );
  NAND3X1 U797 ( .IN1(n686), .IN2(n685), .IN3(n684), .OUT(n687) );
  AOI22 U798 ( .IN1(RSTn), .IN2(n687), .IN3(Final_Mantissa_reg[1]), .IN4(n704), 
        .OUT(n688) );
  INVX1 U799 ( .IN(n688), .OUT(n870) );
  AOI22 U800 ( .IN1(Multi_dataout[8]), .IN2(n716), .IN3(Multi_dataout[7]), 
        .IN4(n113), .OUT(n690) );
  AOI22 U801 ( .IN1(Multi_dataout[9]), .IN2(n717), .IN3(Multi_dataout[6]), 
        .IN4(n114), .OUT(n689) );
  AOI22 U802 ( .IN1(Multi_dataout[4]), .IN2(n716), .IN3(Multi_dataout[3]), 
        .IN4(n113), .OUT(n692) );
  AOI22 U803 ( .IN1(Multi_dataout[5]), .IN2(n717), .IN3(Multi_dataout[2]), 
        .IN4(n114), .OUT(n691) );
  AOI22 U804 ( .IN1(n764), .IN2(n761), .IN3(n762), .IN4(n756), .OUT(n702) );
  OAI21 U805 ( .IN1(n693), .IN2(Final_Mantissa_reg[2]), .IN3(n707), .OUT(n695)
         );
  AOI22 U806 ( .IN1(Multi_dataout[9]), .IN2(n714), .IN3(n497), .IN4(Datain1[2]), .OUT(n694) );
  OAI21 U807 ( .IN1(n512), .IN2(n695), .IN3(n694), .OUT(n700) );
  AOI22 U808 ( .IN1(Multi_dataout[1]), .IN2(n717), .IN3(Multi_dataout[0]), 
        .IN4(n716), .OUT(n697) );
  AOI22 U809 ( .IN1(Multi_dataout[10]), .IN2(n745), .IN3(n498), .IN4(
        Datain2[2]), .OUT(n696) );
  OAI21 U810 ( .IN1(n698), .IN2(n697), .IN3(n696), .OUT(n699) );
  NOR2X1 U811 ( .IN1(n700), .IN2(n699), .OUT(n701) );
  AOI22 U812 ( .IN1(RSTn), .IN2(n705), .IN3(Final_Mantissa_reg[2]), .IN4(n704), 
        .OUT(n706) );
  INVX1 U813 ( .IN(n706), .OUT(n869) );
  AOI22 U814 ( .IN1(Multi_dataout[11]), .IN2(n745), .IN3(Datain2[3]), .IN4(
        n498), .OUT(n713) );
  MUX2X1 U815 ( .IN1(n63), .IN2(Final_Mantissa_reg[3]), .S(n707), .OUT(n708)
         );
  AOI22 U816 ( .IN1(n709), .IN2(n708), .IN3(Datain1[3]), .IN4(n497), .OUT(n712) );
  AOI22 U817 ( .IN1(Multi_dataout[2]), .IN2(n717), .IN3(Multi_dataout[0]), 
        .IN4(n113), .OUT(n710) );
  OAI21 U818 ( .IN1(n225), .IN2(n760), .IN3(n710), .OUT(n788) );
  NAND3X1 U819 ( .IN1(n713), .IN2(n712), .IN3(n711), .OUT(n723) );
  AOI21 U820 ( .IN1(n764), .IN2(n717), .IN3(n714), .OUT(n739) );
  AOI22 U821 ( .IN1(Multi_dataout[8]), .IN2(n113), .IN3(Multi_dataout[7]), 
        .IN4(n114), .OUT(n715) );
  OAI21 U822 ( .IN1(n510), .IN2(n760), .IN3(n715), .OUT(n720) );
  AOI22 U823 ( .IN1(Multi_dataout[5]), .IN2(n716), .IN3(Multi_dataout[4]), 
        .IN4(n113), .OUT(n719) );
  AOI22 U824 ( .IN1(Multi_dataout[6]), .IN2(n717), .IN3(Multi_dataout[3]), 
        .IN4(n114), .OUT(n718) );
  AOI22 U825 ( .IN1(n764), .IN2(n720), .IN3(n762), .IN4(n787), .OUT(n721) );
  OAI21 U826 ( .IN1(n739), .IN2(n176), .IN3(n721), .OUT(n722) );
  OAI21 U827 ( .IN1(n723), .IN2(n722), .IN3(RSTn), .OUT(n724) );
  OAI21 U828 ( .IN1(n771), .IN2(n63), .IN3(n724), .OUT(n868) );
  AOI22 U829 ( .IN1(n498), .IN2(Datain2[4]), .IN3(n497), .IN4(Datain1[4]), 
        .OUT(n731) );
  AOI22 U830 ( .IN1(Multi_dataout[12]), .IN2(n745), .IN3(n726), .IN4(n725), 
        .OUT(n730) );
  AOI21 U831 ( .IN1(n728), .IN2(Final_Mantissa_reg[4]), .IN3(n512), .OUT(n727)
         );
  OAI21 U832 ( .IN1(n728), .IN2(Final_Mantissa_reg[4]), .IN3(n727), .OUT(n729)
         );
  NAND3X1 U833 ( .IN1(n731), .IN2(n730), .IN3(n729), .OUT(n737) );
  AOI22 U834 ( .IN1(Multi_dataout[8]), .IN2(n114), .IN3(Multi_dataout[9]), 
        .IN4(n113), .OUT(n732) );
  OAI21 U835 ( .IN1(n176), .IN2(n760), .IN3(n732), .OUT(n734) );
  AOI22 U836 ( .IN1(n764), .IN2(n734), .IN3(n762), .IN4(n733), .OUT(n735) );
  OAI21 U837 ( .IN1(n739), .IN2(n509), .IN3(n735), .OUT(n736) );
  OAI21 U838 ( .IN1(n737), .IN2(n736), .IN3(RSTn), .OUT(n738) );
  OAI21 U839 ( .IN1(n771), .IN2(n68), .IN3(n738), .OUT(n867) );
  INVX1 U840 ( .IN(n739), .OUT(n744) );
  AOI22 U841 ( .IN1(n498), .IN2(Datain2[6]), .IN3(n497), .IN4(Datain1[6]), 
        .OUT(n751) );
  AOI22 U842 ( .IN1(Multi_dataout[14]), .IN2(n745), .IN3(Multi_dataout[13]), 
        .IN4(n744), .OUT(n750) );
  OAI21 U843 ( .IN1(n748), .IN2(Final_Mantissa_reg[6]), .IN3(n747), .OUT(n749)
         );
  NAND3X1 U844 ( .IN1(n751), .IN2(n750), .IN3(n749), .OUT(n769) );
  OAI21 U845 ( .IN1(Multi_dataout[1]), .IN2(n754), .IN3(n752), .OUT(n753) );
  AOI22 U846 ( .IN1(Multi_dataout[10]), .IN2(n114), .IN3(Multi_dataout[11]), 
        .IN4(n113), .OUT(n759) );
  OAI21 U847 ( .IN1(n508), .IN2(n760), .IN3(n759), .OUT(n763) );
  AOI22 U848 ( .IN1(n764), .IN2(n763), .IN3(n762), .IN4(n761), .OUT(n765) );
  OAI21 U849 ( .IN1(n767), .IN2(n766), .IN3(n765), .OUT(n768) );
  OAI21 U850 ( .IN1(n769), .IN2(n768), .IN3(RSTn), .OUT(n770) );
  OAI21 U851 ( .IN1(n771), .IN2(n73), .IN3(n770), .OUT(n865) );
  NOR2X1 U852 ( .IN1(n52), .IN2(n126), .OUT(n775) );
  NAND3X1 U853 ( .IN1(n772), .IN2(n777), .IN3(n512), .OUT(n773) );
  OAI21 U854 ( .IN1(Dataout_valid), .IN2(n773), .IN3(RSTn), .OUT(n774) );
  MUX2X1 U855 ( .IN1(ExcCheck_valid), .IN2(n775), .S(n774), .OUT(n864) );
  NOR2X1 U856 ( .IN1(StateMC[2]), .IN2(n778), .OUT(n780) );
  AOI21 U857 ( .IN1(n780), .IN2(n779), .IN3(n126), .OUT(n832) );
  NOR2X1 U858 ( .IN1(n789), .IN2(n781), .OUT(n786) );
  AOI22 U859 ( .IN1(Multi_dataout[6]), .IN2(n502), .IN3(Multi_dataout[5]), 
        .IN4(n786), .OUT(n785) );
  NOR2X1 U860 ( .IN1(n795), .IN2(n782), .OUT(n790) );
  AOI22 U861 ( .IN1(n790), .IN2(n783), .IN3(T_reg), .IN4(n789), .OUT(n784) );
  AOI22 U862 ( .IN1(Multi_dataout[7]), .IN2(n502), .IN3(Multi_dataout[6]), 
        .IN4(n786), .OUT(n793) );
  AOI22 U863 ( .IN1(n791), .IN2(n790), .IN3(G_reg), .IN4(n789), .OUT(n792) );
  AOI21 U864 ( .IN1(n474), .IN2(n795), .IN3(n836), .OUT(n796) );
  OAI21 U865 ( .IN1(n796), .IN2(n854), .IN3(n489), .OUT(n828) );
  AOI22 U866 ( .IN1(RSTn), .IN2(n797), .IN3(Debug_reg[1]), .IN4(n828), .OUT(
        n798) );
  OAI21 U867 ( .IN1(n505), .IN2(n853), .IN3(n884), .OUT(n799) );
  NOR2X1 U868 ( .IN1(n833), .IN2(n799), .OUT(n803) );
  OAI21 U869 ( .IN1(n126), .IN2(n836), .IN3(n800), .OUT(n802) );
  AOI22 U870 ( .IN1(Op1_Mantissa_reg[7]), .IN2(n803), .IN3(Multi_datain1[7]), 
        .IN4(n802), .OUT(n801) );
  AOI22 U871 ( .IN1(n803), .IN2(Op1_Mantissa_reg[6]), .IN3(Multi_datain1[6]), 
        .IN4(n802), .OUT(n804) );
  AOI22 U872 ( .IN1(n491), .IN2(Datain2[6]), .IN3(Op2_Mantissa_reg[6]), .IN4(
        n112), .OUT(n805) );
  AOI22 U873 ( .IN1(n491), .IN2(Datain2[5]), .IN3(Op2_Mantissa_reg[5]), .IN4(
        n112), .OUT(n806) );
  AOI22 U874 ( .IN1(n491), .IN2(Datain2[4]), .IN3(Op2_Mantissa_reg[4]), .IN4(
        n112), .OUT(n807) );
  AOI22 U875 ( .IN1(n491), .IN2(Datain2[3]), .IN3(Op2_Mantissa_reg[3]), .IN4(
        n112), .OUT(n808) );
  AOI22 U876 ( .IN1(n491), .IN2(Datain2[2]), .IN3(Op2_Mantissa_reg[2]), .IN4(
        n112), .OUT(n809) );
  AOI22 U877 ( .IN1(n491), .IN2(Datain2[1]), .IN3(Op2_Mantissa_reg[1]), .IN4(
        n112), .OUT(n810) );
  AOI22 U878 ( .IN1(n491), .IN2(Datain2[0]), .IN3(Op2_Mantissa_reg[0]), .IN4(
        n112), .OUT(n811) );
  AOI22 U879 ( .IN1(n491), .IN2(n127), .IN3(Op1_Mantissa_reg[7]), .IN4(n112), 
        .OUT(n812) );
  AOI22 U880 ( .IN1(n491), .IN2(Datain1[6]), .IN3(Op1_Mantissa_reg[6]), .IN4(
        n112), .OUT(n813) );
  AOI22 U881 ( .IN1(n491), .IN2(Datain1[5]), .IN3(Op1_Mantissa_reg[5]), .IN4(
        n112), .OUT(n814) );
  AOI22 U882 ( .IN1(n491), .IN2(Datain1[4]), .IN3(Op1_Mantissa_reg[4]), .IN4(
        n112), .OUT(n815) );
  AOI22 U883 ( .IN1(n491), .IN2(Datain1[3]), .IN3(Op1_Mantissa_reg[3]), .IN4(
        n112), .OUT(n816) );
  AOI22 U884 ( .IN1(n491), .IN2(Datain1[2]), .IN3(Op1_Mantissa_reg[2]), .IN4(
        n112), .OUT(n817) );
  AOI22 U885 ( .IN1(n491), .IN2(Datain1[1]), .IN3(Op1_Mantissa_reg[1]), .IN4(
        n112), .OUT(n818) );
  AOI22 U886 ( .IN1(n491), .IN2(Datain1[0]), .IN3(Op1_Mantissa_reg[0]), .IN4(
        n112), .OUT(n820) );
  NAND3X1 U887 ( .IN1(n499), .IN2(n821), .IN3(n474), .OUT(n826) );
  NAND3X1 U888 ( .IN1(n490), .IN2(Multi_dataout[15]), .IN3(Multi_ack), .OUT(
        n822) );
  OAI21 U889 ( .IN1(n823), .IN2(n826), .IN3(n822), .OUT(n824) );
  AOI22 U890 ( .IN1(n319), .IN2(n824), .IN3(Debug_reg[3]), .IN4(n828), .OUT(
        n825) );
  NOR2X1 U891 ( .IN1(n827), .IN2(n826), .OUT(n829) );
  AOI22 U892 ( .IN1(n319), .IN2(n829), .IN3(Debug_reg[2]), .IN4(n828), .OUT(
        n831) );
  NOR2X1 U893 ( .IN1(n836), .IN2(n854), .OUT(n858) );
  NAND3X1 U894 ( .IN1(n490), .IN2(n858), .IN3(Multi_dataout[14]), .OUT(n830)
         );
  NOR2X1 U895 ( .IN1(n832), .IN2(n491), .OUT(n835) );
  INVX1 U896 ( .IN(n835), .OUT(n834) );
  AOI22 U897 ( .IN1(n835), .IN2(n833), .IN3(Multi_valid_BAR), .IN4(n834), 
        .OUT(n142) );
  NOR2X1 U898 ( .IN1(n834), .IN2(n833), .OUT(n851) );
  OAI21 U899 ( .IN1(n126), .IN2(n836), .IN3(n835), .OUT(n850) );
  AOI22 U900 ( .IN1(Op2_Mantissa_reg[7]), .IN2(n115), .IN3(Multi_datain2[7]), 
        .IN4(n850), .OUT(n837) );
  AOI22 U901 ( .IN1(Op2_Mantissa_reg[6]), .IN2(n115), .IN3(Multi_datain2[6]), 
        .IN4(n850), .OUT(n838) );
  AOI22 U902 ( .IN1(Op2_Mantissa_reg[5]), .IN2(n115), .IN3(Multi_datain2[5]), 
        .IN4(n850), .OUT(n839) );
  AOI22 U903 ( .IN1(Op2_Mantissa_reg[4]), .IN2(n115), .IN3(Multi_datain2[4]), 
        .IN4(n850), .OUT(n840) );
  AOI22 U904 ( .IN1(Op2_Mantissa_reg[3]), .IN2(n115), .IN3(Multi_datain2[3]), 
        .IN4(n850), .OUT(n841) );
  AOI22 U905 ( .IN1(Op2_Mantissa_reg[2]), .IN2(n115), .IN3(Multi_datain2[2]), 
        .IN4(n850), .OUT(n842) );
  AOI22 U906 ( .IN1(Op2_Mantissa_reg[1]), .IN2(n115), .IN3(Multi_datain2[1]), 
        .IN4(n850), .OUT(n843) );
  AOI22 U907 ( .IN1(Op2_Mantissa_reg[0]), .IN2(n115), .IN3(Multi_datain2[0]), 
        .IN4(n850), .OUT(n844) );
  AOI22 U908 ( .IN1(Op1_Mantissa_reg[5]), .IN2(n115), .IN3(Multi_datain1[5]), 
        .IN4(n850), .OUT(n845) );
  AOI22 U909 ( .IN1(Op1_Mantissa_reg[4]), .IN2(n115), .IN3(Multi_datain1[4]), 
        .IN4(n850), .OUT(n846) );
  AOI22 U910 ( .IN1(Op1_Mantissa_reg[3]), .IN2(n115), .IN3(Multi_datain1[3]), 
        .IN4(n850), .OUT(n847) );
  AOI22 U911 ( .IN1(Op1_Mantissa_reg[2]), .IN2(n115), .IN3(Multi_datain1[2]), 
        .IN4(n850), .OUT(n848) );
  AOI22 U912 ( .IN1(Op1_Mantissa_reg[1]), .IN2(n115), .IN3(Multi_datain1[1]), 
        .IN4(n850), .OUT(n849) );
  AOI22 U913 ( .IN1(Op1_Mantissa_reg[0]), .IN2(n115), .IN3(Multi_datain1[0]), 
        .IN4(n850), .OUT(n852) );
  OAI21 U914 ( .IN1(Multi_ack), .IN2(n854), .IN3(n853), .OUT(n859) );
  AOI22 U915 ( .IN1(G_reg), .IN2(n859), .IN3(n858), .IN4(n855), .OUT(n856) );
  INVX1 U916 ( .IN(n856), .OUT(n125) );
  AOI22 U917 ( .IN1(T_reg), .IN2(n859), .IN3(n858), .IN4(n857), .OUT(n860) );
  INVX1 U918 ( .IN(n860), .OUT(n124) );
endmodule


module FPU_Control ( CLK, RSTn, CS, DIN1, DIN2, DIV, DACK, DR, DOUT, DOV, DOA, 
        ABUSY, MBUSY, EXC, OPT, MODE, DEBUG );
  input [15:0] DIN1;
  input [15:0] DIN2;
  output [15:0] DOUT;
  output [2:0] EXC;
  input [2:0] MODE;
  output [4:0] DEBUG;
  input CLK, RSTn, CS, DIV, DOA, OPT;
  output DACK, DR, DOV, ABUSY, MBUSY;
  wire   Add_carryout, N149, N150, N151, N152, N191, N192, N193,
         MulCntrl_valid, AdderCntrl_valid, AdderCntrl_Dataout_valid,
         MulCntrl_Dataout_valid, Add_valid, Add_ack, AdderCntrl_ExcCheck_valid,
         AdderCntrl_Exc_Ack, Booth_valid, Booth_ack, MulCntrl_ExcCheck_valid,
         MulCntrl_Exc_Ack, ExcSelect, ExcCheck_valid, Booth_Add_valid,
         Booth_Add_ack, AddSelect, u_exc_check_N45, u_exc_check_StateMC_0_,
         u_ExcChecker_interconnect_N53, u_ExcChecker_interconnect_priority_reg,
         u_ExcChecker_interconnect_stateMC_0_,
         u_ExcChecker_interconnect_stateMC_1_, u_booth_N258, u_booth_N55,
         u_booth_N54, u_booth_N53, u_booth_N52, u_booth_N51, u_booth_N50,
         u_booth_N49, u_booth_BStateMC_1_, u_booth_count_reg_2_,
         u_booth_count_reg_3_, u_booth_Q1_reg, u_booth_M_reg_1_,
         u_booth_M_reg_2_, u_booth_M_reg_3_, u_booth_M_reg_4_,
         u_booth_M_reg_5_, u_booth_M_reg_6_, u_booth_M_reg_7_,
         u_booth_A_reg_7_, u_booth_A_reg_8_, u_adder_24b_N131,
         u_adder_24b_N130, u_adder_24b_N129, u_adder_24b_N128,
         u_adder_24b_N127, u_adder_24b_N126, u_adder_24b_N125,
         u_adder_24b_N124, u_adder_24b_N123, u_adder_24b_N122, u_adder_24b_N52,
         u_adder_24b_StateMC_1_, u_Adder_interconnect_N53,
         u_Adder_interconnect_priority_reg, u_Adder_interconnect_stateMC_1_,
         n408, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n462, n463,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n587, n588, n592, n594,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n610,
         n611, n612, n613, n614, n615, n616, n617, n622, n654, n694, n695,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n732, n768, n802, n806, n992, n1022,
         n1028, n1031, n1034, n1037, n1040, n1043, n1077, n1079, n1088, n1092,
         n1135, n1302, n1513, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1587, n1588, n1589, n1620,
         n1621, n1622, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1692, n1723, add_x_176_n13, add_x_176_n12, add_x_176_n11,
         add_x_176_n10, add_x_176_n9, add_x_176_n8, add_x_176_n7, add_x_176_n6,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2;
  wire   [8:0] Add_dataout;
  wire   [4:0] AdderCntrl_Debug;
  wire   [1:0] multStateMC;
  wire   [4:0] MulCntrl_Debug;
  wire   [15:0] AdderCntrl_Op1;
  wire   [15:0] AdderCntrl_Op2;
  wire   [15:0] MulCntrl_Op1;
  wire   [15:0] MulCntrl_Op2;
  wire   [1:0] getdataStat_reg;
  wire   [15:0] AdderResult_reg;
  wire   [15:0] MultResult_reg;
  wire   [2:0] AddExc_reg;
  wire   [2:0] MultExc_reg;
  wire   [15:0] AdderCntrl_Dataout;
  wire   [2:0] AdderCntrl_Exc;
  wire   [15:0] MulCntrl_Dataout;
  wire   [2:0] MulCntrl_Exc;
  wire   [7:0] Add_Op1;
  wire   [8:0] Add_Op2;
  wire   [14:0] AdderCntrl_ExcCheck_Datain;
  wire   [2:0] ExcCheck_value;
  wire   [7:0] Booth_datain1;
  wire   [7:0] Booth_datain2;
  wire   [15:0] Booth_dataout;
  wire   [14:0] MulCntrl_ExcCheck_Datain;
  wire   [8:0] Booth_Add_datain1;
  wire   [8:0] Booth_Add_datain2;
  wire   [8:0] Add_Op1_wire;
  wire   [8:1] Add_Op2_wire;

  Adder_cntrl u_adder_cntrl ( .CLK(CLK), .RSTn(n1794), .Datain1(AdderCntrl_Op1), .Datain2(AdderCntrl_Op2), .Data_valid(AdderCntrl_valid), .Dataout(
        AdderCntrl_Dataout), .Exc(AdderCntrl_Exc), .Mode(MODE), .Debug(
        AdderCntrl_Debug), .Adder_datain1({SYNOPSYS_UNCONNECTED_1, Add_Op1}), 
        .Adder_datain2(Add_Op2), .Adder_valid(Add_valid), .Adder_dataout(
        Add_dataout), .Adder_carryout(Add_carryout), .Adder_ack(Add_ack), 
        .ExcCheck_valid(AdderCntrl_ExcCheck_valid), .Exc_value(ExcCheck_value), 
        .Exc_Ack(AdderCntrl_Exc_Ack), .Dataout_valid_BAR(
        AdderCntrl_Dataout_valid), .ExcCheck_Datain_14_(
        AdderCntrl_ExcCheck_Datain[14]), .ExcCheck_Datain_13__BAR(
        AdderCntrl_ExcCheck_Datain[13]), .ExcCheck_Datain_12_(
        AdderCntrl_ExcCheck_Datain[12]), .ExcCheck_Datain_11_(
        AdderCntrl_ExcCheck_Datain[11]), .ExcCheck_Datain_9_(
        AdderCntrl_ExcCheck_Datain[9]), .ExcCheck_Datain_8_(
        AdderCntrl_ExcCheck_Datain[8]), .ExcCheck_Datain_6_(
        AdderCntrl_ExcCheck_Datain[6]), .ExcCheck_Datain_5_(
        AdderCntrl_ExcCheck_Datain[5]), .ExcCheck_Datain_4_(
        AdderCntrl_ExcCheck_Datain[4]), .ExcCheck_Datain_3_(
        AdderCntrl_ExcCheck_Datain[3]), .ExcCheck_Datain_2_(
        AdderCntrl_ExcCheck_Datain[2]), .ExcCheck_Datain_1_(
        AdderCntrl_ExcCheck_Datain[1]), .ExcCheck_Datain_0_(
        AdderCntrl_ExcCheck_Datain[0]), .ExcCheck_Datain_10__BAR(
        AdderCntrl_ExcCheck_Datain[10]), .ExcCheck_Datain_7__BAR(
        AdderCntrl_ExcCheck_Datain[7]) );
  Mul_cntrl u_mul_cntrl ( .CLK(CLK), .RSTn(n1794), .Datain1({
        MulCntrl_Op1[15:8], n1733, MulCntrl_Op1[6:0]}), .Datain2({
        MulCntrl_Op2[15:8], n1735, MulCntrl_Op2[6:0]}), .Data_valid(
        MulCntrl_valid), .Dataout(MulCntrl_Dataout), .Dataout_valid(
        MulCntrl_Dataout_valid), .Exc(MulCntrl_Exc), .Mode(MODE), .Debug(
        MulCntrl_Debug), .Multi_datain1(Booth_datain1), .Multi_datain2(
        Booth_datain2), .Multi_dataout(Booth_dataout), .Multi_ack(Booth_ack), 
        .ExcCheck_valid(MulCntrl_ExcCheck_valid), .ExcCheck_Datain({
        SYNOPSYS_UNCONNECTED_2, MulCntrl_ExcCheck_Datain}), .Exc_value(
        ExcCheck_value), .Multi_valid_BAR(Booth_valid), .Exc_Ack_BAR(n1730) );
  DFFRX1 u_Adder_interconnect_M2_ack_reg ( .D(n1587), .CLK(CLK), .CLRB(n408), 
        .Q(Booth_Add_ack), .QB(n1745) );
  DFFRX1 u_booth_count_reg_reg_0_ ( .D(n1554), .CLK(CLK), .CLRB(n408), .QB(
        n694) );
  DFFRX1 u_booth_count_reg_reg_1_ ( .D(n1079), .CLK(CLK), .CLRB(n408), .Q(n695) );
  DFFRX1 u_booth_count_reg_reg_2_ ( .D(n1555), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_count_reg_2_) );
  DFFRX1 u_booth_count_reg_reg_3_ ( .D(n1092), .CLK(CLK), .CLRB(n408), .Q(
        n1767), .QB(u_booth_count_reg_3_) );
  DFFRX1 u_booth_BStateMC_reg_0_ ( .D(n1556), .CLK(CLK), .CLRB(n408), .Q(n1781), .QB(n732) );
  DFFRX1 u_booth_BStateMC_reg_1_ ( .D(n1088), .CLK(CLK), .CLRB(n408), .Q(n1780), .QB(u_booth_BStateMC_1_) );
  DFFRX1 u_booth_Q_reg_reg_7_ ( .D(n1022), .CLK(CLK), .CLRB(n408), .Q(n720), 
        .QB(n1759) );
  DFFRX1 u_booth_Q_reg_reg_6_ ( .D(n1028), .CLK(CLK), .CLRB(n408), .Q(n719), 
        .QB(n1760) );
  DFFRX1 u_booth_Q_reg_reg_5_ ( .D(n1031), .CLK(CLK), .CLRB(n408), .Q(n718), 
        .QB(n1761) );
  DFFRX1 u_booth_Q_reg_reg_4_ ( .D(n1034), .CLK(CLK), .CLRB(n408), .Q(n717), 
        .QB(n1762) );
  DFFRX1 u_booth_Q_reg_reg_3_ ( .D(n1037), .CLK(CLK), .CLRB(n408), .Q(n716), 
        .QB(n1763) );
  DFFRX1 u_booth_Q_reg_reg_2_ ( .D(n1040), .CLK(CLK), .CLRB(n408), .Q(n715), 
        .QB(n1764) );
  DFFRX1 u_booth_Q_reg_reg_1_ ( .D(n1043), .CLK(CLK), .CLRB(n408), .Q(n714), 
        .QB(n1765) );
  DFFRX1 u_booth_Q_reg_reg_0_ ( .D(n1135), .CLK(CLK), .CLRB(n408), .Q(n713), 
        .QB(n1736) );
  DFFRX1 u_booth_Adder_valid_reg ( .D(n1653), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_valid), .QB(n1758) );
  DFFRX1 u_Adder_interconnect_priority_reg_reg ( .D(n1620), .CLK(CLK), .CLRB(
        n408), .Q(u_Adder_interconnect_priority_reg), .QB(n1740) );
  DFFRX1 u_Adder_interconnect_stateMC_reg_0_ ( .D(n1621), .CLK(CLK), .CLRB(
        n408), .Q(n1739), .QB(n806) );
  DFFRX1 u_Adder_interconnect_M1_ack_reg ( .D(n594), .CLK(CLK), .CLRB(n408), 
        .Q(Add_ack) );
  DFFRX1 u_ExcChecker_interconnect_stateMC_reg_1_ ( .D(n1661), .CLK(CLK), 
        .CLRB(n408), .Q(u_ExcChecker_interconnect_stateMC_1_), .QB(n1755) );
  DFFRX1 u_ExcChecker_interconnect_priority_reg_reg ( .D(n1659), .CLK(CLK), 
        .CLRB(n408), .Q(u_ExcChecker_interconnect_priority_reg), .QB(n1752) );
  DFFRX1 u_ExcChecker_interconnect_stateMC_reg_0_ ( .D(n1660), .CLK(CLK), 
        .CLRB(n408), .Q(u_ExcChecker_interconnect_stateMC_0_), .QB(n1753) );
  DFFRX1 u_ExcChecker_interconnect_S_req_reg ( .D(
        u_ExcChecker_interconnect_N53), .CLK(CLK), .CLRB(n408), .Q(
        ExcCheck_valid) );
  DFFRX1 u_exc_check_ACK_reg ( .D(u_exc_check_N45), .CLK(CLK), .CLRB(n408), 
        .QB(n1748) );
  DFFRX1 u_ExcChecker_interconnect_M2_ack_reg ( .D(n1656), .CLK(CLK), .CLRB(
        n408), .Q(MulCntrl_Exc_Ack), .QB(n1730) );
  DFFRX1 u_exc_check_StateMC_reg_0_ ( .D(n622), .CLK(CLK), .CLRB(n408), .Q(
        u_exc_check_StateMC_0_), .QB(n1766) );
  DFFRX1 u_exc_check_StateMC_reg_1_ ( .D(n1657), .CLK(CLK), .CLRB(n408), .Q(
        n1772), .QB(n654) );
  DFFRX1 u_ExcChecker_interconnect_Select_reg ( .D(n1658), .CLK(CLK), .CLRB(
        n408), .Q(ExcSelect), .QB(n1747) );
  DFFRX1 u_exc_check_AEXC_reg_2_ ( .D(n588), .CLK(CLK), .CLRB(n408), .Q(
        ExcCheck_value[2]) );
  DFFRX1 u_exc_check_AEXC_reg_1_ ( .D(n1654), .CLK(CLK), .CLRB(n408), .Q(
        ExcCheck_value[1]), .QB(n1751) );
  DFFRX1 u_exc_check_AEXC_reg_0_ ( .D(n1655), .CLK(CLK), .CLRB(n408), .Q(
        ExcCheck_value[0]), .QB(n1769) );
  DFFRX1 u_ExcChecker_interconnect_M1_ack_reg ( .D(n592), .CLK(CLK), .CLRB(
        n408), .Q(AdderCntrl_Exc_Ack) );
  DFFRX1 u_Adder_interconnect_stateMC_reg_1_ ( .D(n1622), .CLK(CLK), .CLRB(
        n408), .Q(u_Adder_interconnect_stateMC_1_), .QB(n1754) );
  DFFRX1 u_Adder_interconnect_S_req_reg ( .D(u_Adder_interconnect_N53), .CLK(
        CLK), .CLRB(n408), .QB(n802) );
  DFFRX1 u_adder_24b_StateMC_reg_1_ ( .D(n1589), .CLK(CLK), .CLRB(n408), .Q(
        u_adder_24b_StateMC_1_), .QB(n1757) );
  DFFRX1 u_adder_24b_StateMC_reg_0_ ( .D(n1588), .CLK(CLK), .CLRB(n408), .Q(
        n1770), .QB(n768) );
  DFFRX1 u_adder_24b_ACK_reg ( .D(u_adder_24b_N52), .CLK(CLK), .CLRB(n408), 
        .QB(n1749) );
  DFFRX1 u_adder_24b_Z_reg_8_ ( .D(n598), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[8]) );
  DFFRX1 u_adder_24b_Z_reg_7_ ( .D(n599), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[7]) );
  DFFRX1 u_adder_24b_Z_reg_6_ ( .D(n600), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[6]) );
  DFFRX1 u_adder_24b_Z_reg_5_ ( .D(n601), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[5]) );
  DFFRX1 u_adder_24b_Z_reg_4_ ( .D(n602), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[4]) );
  DFFRX1 u_adder_24b_Z_reg_3_ ( .D(n603), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[3]) );
  DFFRX1 u_adder_24b_Z_reg_2_ ( .D(n604), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[2]) );
  DFFRX1 u_adder_24b_Z_reg_1_ ( .D(n605), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[1]) );
  DFFRX1 u_adder_24b_Z_reg_0_ ( .D(n596), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[0]) );
  DFFRX1 u_adder_24b_COUT_reg ( .D(n597), .CLK(CLK), .CLRB(n408), .Q(
        Add_carryout) );
  DFFRX1 adderStateMC_reg_0_ ( .D(n1302), .CLK(CLK), .CLRB(n408), .Q(n463), 
        .QB(n1744) );
  DFFRX1 outputRdy_reg_reg_0_ ( .D(N191), .CLK(CLK), .CLRB(n408), .QB(n587) );
  DFFRX1 adderStateMC_reg_1_ ( .D(n1692), .CLK(CLK), .CLRB(n408), .Q(n1741), 
        .QB(n462) );
  DFFRX1 getdataStat_reg_reg_0_ ( .D(N149), .CLK(CLK), .CLRB(n408), .Q(
        getdataStat_reg[0]) );
  DFFRX1 AdderCntrl_Op2_reg_0_ ( .D(n551), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[0]) );
  DFFRX1 AdderCntrl_Op2_reg_1_ ( .D(n550), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[1]) );
  DFFRX1 AdderCntrl_Op2_reg_2_ ( .D(n549), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[2]) );
  DFFRX1 AdderCntrl_Op2_reg_3_ ( .D(n548), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[3]) );
  DFFRX1 AdderCntrl_Op2_reg_4_ ( .D(n547), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[4]) );
  DFFRX1 AdderCntrl_Op2_reg_5_ ( .D(n546), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[5]) );
  DFFRX1 AdderCntrl_Op2_reg_6_ ( .D(n545), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[6]) );
  DFFRX1 AdderCntrl_Op2_reg_7_ ( .D(n544), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[7]) );
  DFFRX1 AdderCntrl_Op2_reg_8_ ( .D(n543), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[8]) );
  DFFRX1 AdderCntrl_Op2_reg_9_ ( .D(n542), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[9]) );
  DFFRX1 AdderCntrl_Op2_reg_10_ ( .D(n541), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[10]) );
  DFFRX1 AdderCntrl_Op2_reg_11_ ( .D(n540), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[11]) );
  DFFRX1 AdderCntrl_Op2_reg_12_ ( .D(n539), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[12]) );
  DFFRX1 AdderCntrl_Op2_reg_13_ ( .D(n538), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[13]) );
  DFFRX1 AdderCntrl_Op2_reg_14_ ( .D(n537), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[14]) );
  DFFRX1 AdderCntrl_Op2_reg_15_ ( .D(n536), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[15]) );
  DFFRX1 AdderCntrl_Op1_reg_0_ ( .D(n535), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[0]) );
  DFFRX1 AdderCntrl_Op1_reg_1_ ( .D(n534), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[1]) );
  DFFRX1 AdderCntrl_Op1_reg_2_ ( .D(n533), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[2]) );
  DFFRX1 AdderCntrl_Op1_reg_3_ ( .D(n532), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[3]) );
  DFFRX1 AdderCntrl_Op1_reg_4_ ( .D(n531), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[4]) );
  DFFRX1 AdderCntrl_Op1_reg_5_ ( .D(n530), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[5]) );
  DFFRX1 AdderCntrl_Op1_reg_6_ ( .D(n529), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[6]) );
  DFFRX1 AdderCntrl_Op1_reg_7_ ( .D(n528), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[7]) );
  DFFRX1 AdderCntrl_Op1_reg_8_ ( .D(n527), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[8]) );
  DFFRX1 AdderCntrl_Op1_reg_9_ ( .D(n526), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[9]) );
  DFFRX1 AdderCntrl_Op1_reg_10_ ( .D(n525), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[10]) );
  DFFRX1 AdderCntrl_Op1_reg_11_ ( .D(n524), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[11]) );
  DFFRX1 AdderCntrl_Op1_reg_12_ ( .D(n523), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[12]) );
  DFFRX1 AdderCntrl_Op1_reg_13_ ( .D(n522), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[13]) );
  DFFRX1 AdderCntrl_Op1_reg_14_ ( .D(n521), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[14]) );
  DFFRX1 AdderCntrl_Op1_reg_15_ ( .D(n520), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[15]) );
  DFFRX1 ABUSY_reg ( .D(N151), .CLK(CLK), .CLRB(n408), .Q(ABUSY) );
  DFFRX1 AddExc_reg_reg_2_ ( .D(n414), .CLK(CLK), .CLRB(n408), .Q(
        AddExc_reg[2]) );
  DFFRX1 AddExc_reg_reg_1_ ( .D(n413), .CLK(CLK), .CLRB(n408), .Q(
        AddExc_reg[1]) );
  DFFRX1 AddExc_reg_reg_0_ ( .D(n412), .CLK(CLK), .CLRB(n408), .Q(
        AddExc_reg[0]) );
  DFFRX1 AdderResult_reg_reg_0_ ( .D(n415), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[0]) );
  DFFRX1 AdderResult_reg_reg_1_ ( .D(n416), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[1]) );
  DFFRX1 AdderResult_reg_reg_2_ ( .D(n417), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[2]) );
  DFFRX1 AdderResult_reg_reg_3_ ( .D(n418), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[3]) );
  DFFRX1 AdderResult_reg_reg_4_ ( .D(n419), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[4]) );
  DFFRX1 AdderResult_reg_reg_5_ ( .D(n420), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[5]) );
  DFFRX1 AdderResult_reg_reg_6_ ( .D(n421), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[6]) );
  DFFRX1 AdderResult_reg_reg_7_ ( .D(n422), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[7]) );
  DFFRX1 AdderResult_reg_reg_8_ ( .D(n423), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[8]) );
  DFFRX1 AdderResult_reg_reg_9_ ( .D(n424), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[9]) );
  DFFRX1 AdderResult_reg_reg_10_ ( .D(n425), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[10]) );
  DFFRX1 AdderResult_reg_reg_11_ ( .D(n426), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[11]) );
  DFFRX1 AdderResult_reg_reg_12_ ( .D(n427), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[12]) );
  DFFRX1 AdderResult_reg_reg_13_ ( .D(n428), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[13]) );
  DFFRX1 AdderResult_reg_reg_14_ ( .D(n429), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[14]) );
  DFFRX1 AdderResult_reg_reg_15_ ( .D(n430), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[15]) );
  DFFRX1 u_booth_Q1_reg_reg ( .D(n1077), .CLK(CLK), .CLRB(n408), .Q(n1743), 
        .QB(u_booth_Q1_reg) );
  DFFRX1 u_booth_A_reg_reg_8_ ( .D(n1545), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_A_reg_8_), .QB(n1771) );
  DFFRX1 u_booth_A_reg_reg_7_ ( .D(n1546), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_A_reg_7_), .QB(n1756) );
  DFFRX1 u_booth_A_reg_reg_6_ ( .D(n1547), .CLK(CLK), .CLRB(n408), .Q(n1774), 
        .QB(n728) );
  DFFRX1 u_booth_A_reg_reg_5_ ( .D(n1548), .CLK(CLK), .CLRB(n408), .Q(n1773), 
        .QB(n727) );
  DFFRX1 u_booth_A_reg_reg_4_ ( .D(n1549), .CLK(CLK), .CLRB(n408), .Q(n1778), 
        .QB(n726) );
  DFFRX1 u_booth_A_reg_reg_3_ ( .D(n1550), .CLK(CLK), .CLRB(n408), .Q(n1775), 
        .QB(n725) );
  DFFRX1 u_booth_A_reg_reg_2_ ( .D(n1551), .CLK(CLK), .CLRB(n408), .Q(n1776), 
        .QB(n724) );
  DFFRX1 u_booth_A_reg_reg_1_ ( .D(n1552), .CLK(CLK), .CLRB(n408), .Q(n1777), 
        .QB(n723) );
  DFFRX1 u_booth_A_reg_reg_0_ ( .D(n1553), .CLK(CLK), .CLRB(n408), .Q(n1779), 
        .QB(n722) );
  DFFRX1 u_booth_Adder_datain1_reg_0_ ( .D(u_booth_N49), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[0]) );
  DFFRX1 u_booth_Q_reg_reg_8_ ( .D(n1544), .CLK(CLK), .CLRB(n408), .Q(n1768), 
        .QB(n721) );
  DFFRX1 u_booth_Adder_datain1_reg_1_ ( .D(u_booth_N50), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[1]) );
  DFFRX1 u_booth_Adder_datain1_reg_2_ ( .D(u_booth_N51), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[2]) );
  DFFRX1 u_booth_Adder_datain1_reg_3_ ( .D(u_booth_N52), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[3]) );
  DFFRX1 u_booth_Adder_datain1_reg_4_ ( .D(u_booth_N53), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[4]) );
  DFFRX1 u_booth_Adder_datain1_reg_5_ ( .D(u_booth_N54), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[5]) );
  DFFRX1 u_booth_Adder_datain1_reg_6_ ( .D(u_booth_N55), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[6]) );
  DFFRX1 u_booth_Adder_datain1_reg_7_ ( .D(n706), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain1[7]) );
  DFFRX1 u_booth_Adder_datain1_reg_8_ ( .D(n707), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain1[8]) );
  DFFRX1 u_booth_Adder_datain2_reg_8_ ( .D(n705), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[8]) );
  DFFRX1 u_booth_M_reg_reg_0_ ( .D(n610), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_N258), .QB(n1737) );
  DFFRX1 u_booth_Adder_datain2_reg_0_ ( .D(n697), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[0]) );
  DFFRX1 u_booth_M_reg_reg_1_ ( .D(n611), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_1_), .QB(n1742) );
  DFFRX1 u_booth_Adder_datain2_reg_1_ ( .D(n698), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[1]) );
  DFFRX1 u_booth_M_reg_reg_2_ ( .D(n612), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_2_) );
  DFFRX1 u_booth_Adder_datain2_reg_2_ ( .D(n699), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[2]) );
  DFFRX1 u_booth_M_reg_reg_3_ ( .D(n613), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_3_) );
  DFFRX1 u_booth_Adder_datain2_reg_3_ ( .D(n700), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[3]) );
  DFFRX1 u_booth_M_reg_reg_4_ ( .D(n614), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_4_) );
  DFFRX1 u_booth_Adder_datain2_reg_4_ ( .D(n701), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[4]) );
  DFFRX1 u_booth_M_reg_reg_5_ ( .D(n615), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_5_) );
  DFFRX1 u_booth_Adder_datain2_reg_5_ ( .D(n702), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[5]) );
  DFFRX1 u_booth_M_reg_reg_6_ ( .D(n616), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_6_) );
  DFFRX1 u_booth_Adder_datain2_reg_6_ ( .D(n703), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[6]) );
  DFFRX1 u_booth_M_reg_reg_7_ ( .D(n617), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_7_), .QB(n1750) );
  DFFRX1 u_booth_Adder_datain2_reg_7_ ( .D(n704), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[7]) );
  DFFRX1 multStateMC_reg_0_ ( .D(n992), .CLK(CLK), .CLRB(n408), .Q(n1746), 
        .QB(multStateMC[0]) );
  DFFRX1 outputRdy_reg_reg_1_ ( .D(N192), .CLK(CLK), .CLRB(n408), .QB(n584) );
  DFFRX1 multStateMC_reg_1_ ( .D(n1513), .CLK(CLK), .CLRB(n408), .Q(
        multStateMC[1]), .QB(n1738) );
  DFFRX1 getdataStat_reg_reg_1_ ( .D(N150), .CLK(CLK), .CLRB(n408), .Q(
        getdataStat_reg[1]) );
  DFFRX1 MulCntrl_Op2_reg_0_ ( .D(n583), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[0]) );
  DFFRX1 MulCntrl_Op2_reg_1_ ( .D(n582), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[1]) );
  DFFRX1 MulCntrl_Op2_reg_2_ ( .D(n581), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[2]) );
  DFFRX1 MulCntrl_Op2_reg_3_ ( .D(n580), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[3]) );
  DFFRX1 MulCntrl_Op2_reg_4_ ( .D(n579), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[4]) );
  DFFRX1 MulCntrl_Op2_reg_5_ ( .D(n578), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[5]) );
  DFFRX1 MulCntrl_Op2_reg_6_ ( .D(n577), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[6]) );
  DFFRX1 MulCntrl_Op2_reg_7_ ( .D(n576), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[7]), .QB(n1734) );
  DFFRX1 MulCntrl_Op2_reg_8_ ( .D(n575), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[8]) );
  DFFRX1 MulCntrl_Op2_reg_9_ ( .D(n574), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[9]) );
  DFFRX1 MulCntrl_Op2_reg_10_ ( .D(n573), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[10]) );
  DFFRX1 MulCntrl_Op2_reg_11_ ( .D(n572), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[11]) );
  DFFRX1 MulCntrl_Op2_reg_12_ ( .D(n571), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[12]) );
  DFFRX1 MulCntrl_Op2_reg_13_ ( .D(n570), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[13]) );
  DFFRX1 MulCntrl_Op2_reg_14_ ( .D(n569), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[14]) );
  DFFRX1 MulCntrl_Op2_reg_15_ ( .D(n568), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[15]) );
  DFFRX1 MulCntrl_Op1_reg_0_ ( .D(n567), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[0]) );
  DFFRX1 MulCntrl_Op1_reg_1_ ( .D(n566), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[1]) );
  DFFRX1 MulCntrl_Op1_reg_2_ ( .D(n565), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[2]) );
  DFFRX1 MulCntrl_Op1_reg_3_ ( .D(n564), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[3]) );
  DFFRX1 MulCntrl_Op1_reg_4_ ( .D(n563), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[4]) );
  DFFRX1 MulCntrl_Op1_reg_5_ ( .D(n562), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[5]) );
  DFFRX1 MulCntrl_Op1_reg_6_ ( .D(n561), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[6]) );
  DFFRX1 MulCntrl_Op1_reg_7_ ( .D(n560), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[7]) );
  DFFRX1 MulCntrl_Op1_reg_8_ ( .D(n559), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[8]) );
  DFFRX1 MulCntrl_Op1_reg_9_ ( .D(n558), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[9]) );
  DFFRX1 MulCntrl_Op1_reg_10_ ( .D(n557), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[10]) );
  DFFRX1 MulCntrl_Op1_reg_11_ ( .D(n556), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[11]) );
  DFFRX1 MulCntrl_Op1_reg_12_ ( .D(n555), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[12]) );
  DFFRX1 MulCntrl_Op1_reg_13_ ( .D(n554), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[13]) );
  DFFRX1 MulCntrl_Op1_reg_14_ ( .D(n553), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[14]) );
  DFFRX1 MulCntrl_Op1_reg_15_ ( .D(n552), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[15]) );
  DFFRX1 MBUSY_reg ( .D(N152), .CLK(CLK), .CLRB(n408), .Q(MBUSY) );
  DFFRX1 DR_reg ( .D(N193), .CLK(CLK), .CLRB(n408), .Q(DR) );
  DFFRX1 MultExc_reg_reg_2_ ( .D(n469), .CLK(CLK), .CLRB(n408), .Q(
        MultExc_reg[2]) );
  DFFRX1 MultExc_reg_reg_1_ ( .D(n468), .CLK(CLK), .CLRB(n408), .Q(
        MultExc_reg[1]) );
  DFFRX1 MultExc_reg_reg_0_ ( .D(n467), .CLK(CLK), .CLRB(n408), .Q(
        MultExc_reg[0]) );
  DFFRX1 MultResult_reg_reg_0_ ( .D(n470), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[0]) );
  DFFRX1 MultResult_reg_reg_1_ ( .D(n471), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[1]) );
  DFFRX1 MultResult_reg_reg_2_ ( .D(n472), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[2]) );
  DFFRX1 MultResult_reg_reg_3_ ( .D(n473), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[3]) );
  DFFRX1 MultResult_reg_reg_4_ ( .D(n474), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[4]) );
  DFFRX1 MultResult_reg_reg_5_ ( .D(n475), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[5]) );
  DFFRX1 MultResult_reg_reg_6_ ( .D(n476), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[6]) );
  DFFRX1 MultResult_reg_reg_7_ ( .D(n477), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[7]) );
  DFFRX1 MultResult_reg_reg_8_ ( .D(n478), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[8]) );
  DFFRX1 MultResult_reg_reg_9_ ( .D(n479), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[9]) );
  DFFRX1 MultResult_reg_reg_10_ ( .D(n480), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[10]) );
  DFFRX1 MultResult_reg_reg_11_ ( .D(n481), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[11]) );
  DFFRX1 MultResult_reg_reg_12_ ( .D(n482), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[12]) );
  DFFRX1 MultResult_reg_reg_13_ ( .D(n483), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[13]) );
  DFFRX1 MultResult_reg_reg_14_ ( .D(n484), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[14]) );
  DFFRX1 MultResult_reg_reg_15_ ( .D(n485), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[15]) );
  DFFRX1 u_Adder_interconnect_Select_reg ( .D(n1723), .CLK(CLK), .CLRB(n408), 
        .Q(AddSelect) );
  FULLADD add_x_176_U9 ( .A(Add_Op1_wire[1]), .B(Add_Op2_wire[1]), .CIN(
        add_x_176_n13), .COUT(add_x_176_n12), .SUM(u_adder_24b_N123) );
  FULLADD add_x_176_U8 ( .A(Add_Op1_wire[2]), .B(Add_Op2_wire[2]), .CIN(
        add_x_176_n12), .COUT(add_x_176_n11), .SUM(u_adder_24b_N124) );
  FULLADD add_x_176_U7 ( .A(Add_Op1_wire[3]), .B(Add_Op2_wire[3]), .CIN(
        add_x_176_n11), .COUT(add_x_176_n10), .SUM(u_adder_24b_N125) );
  FULLADD add_x_176_U6 ( .A(Add_Op1_wire[4]), .B(Add_Op2_wire[4]), .CIN(
        add_x_176_n10), .COUT(add_x_176_n9), .SUM(u_adder_24b_N126) );
  FULLADD add_x_176_U5 ( .A(Add_Op1_wire[5]), .B(Add_Op2_wire[5]), .CIN(
        add_x_176_n9), .COUT(add_x_176_n8), .SUM(u_adder_24b_N127) );
  FULLADD add_x_176_U4 ( .A(Add_Op1_wire[6]), .B(Add_Op2_wire[6]), .CIN(
        add_x_176_n8), .COUT(add_x_176_n7), .SUM(u_adder_24b_N128) );
  FULLADD add_x_176_U3 ( .A(Add_Op1_wire[7]), .B(Add_Op2_wire[7]), .CIN(
        add_x_176_n7), .COUT(add_x_176_n6), .SUM(u_adder_24b_N129) );
  FULLADD add_x_176_U2 ( .A(Add_Op1_wire[8]), .B(Add_Op2_wire[8]), .CIN(
        add_x_176_n6), .COUT(u_adder_24b_N131), .SUM(u_adder_24b_N130) );
  NAND2X1 U1588 ( .IN1(n1780), .IN2(n1781), .OUT(n1725) );
  INVX1 U1589 ( .IN(n1725), .OUT(n1830) );
  NAND3X1 U1590 ( .IN1(n1794), .IN2(Booth_valid), .IN3(n732), .OUT(n1726) );
  NAND2X1 U1591 ( .IN1(n1864), .IN2(n1726), .OUT(n1860) );
  INVX1 U1592 ( .IN(n1830), .OUT(n1727) );
  NOR2X1 U1593 ( .IN1(n2006), .IN2(n1727), .OUT(n1846) );
  NAND3X1 U1594 ( .IN1(n2021), .IN2(n1861), .IN3(Booth_Add_ack), .OUT(n1728)
         );
  INVX1 U1595 ( .IN(n1728), .OUT(n1866) );
  INVX1 U1596 ( .IN(n1853), .OUT(n1729) );
  NOR2X1 U1597 ( .IN1(Booth_valid), .IN2(n1729), .OUT(n1845) );
  INVX4 U1598 ( .IN(AdderCntrl_ExcCheck_Datain[7]), .OUT(n1731) );
  INVX4 U1599 ( .IN(AdderCntrl_ExcCheck_Datain[10]), .OUT(n1732) );
  INVX1 U1600 ( .IN(n2087), .OUT(n601) );
  INVX1 U1601 ( .IN(n2086), .OUT(n602) );
  INVX1 U1602 ( .IN(n2110), .OUT(n588) );
  INVX1 U1603 ( .IN(n2085), .OUT(n603) );
  INVX1 U1604 ( .IN(n2084), .OUT(n604) );
  INVX1 U1605 ( .IN(n2048), .OUT(n703) );
  INVX1 U1606 ( .IN(n2155), .OUT(n543) );
  INVX1 U1607 ( .IN(n2180), .OUT(n520) );
  INVX1 U1608 ( .IN(n2115), .OUT(n580) );
  INVX1 U1609 ( .IN(n2169), .OUT(n529) );
  INVX1 U1610 ( .IN(n2125), .OUT(n570) );
  INVX1 U1611 ( .IN(n2083), .OUT(n605) );
  INVX1 U1612 ( .IN(n2114), .OUT(n581) );
  INVX1 U1613 ( .IN(n2163), .OUT(n535) );
  INVX1 U1614 ( .IN(n2164), .OUT(n534) );
  INVX1 U1615 ( .IN(n2113), .OUT(n582) );
  INVX1 U1616 ( .IN(n2168), .OUT(n530) );
  INVX1 U1617 ( .IN(n2174), .OUT(n524) );
  INVX1 U1618 ( .IN(n2165), .OUT(n533) );
  INVX1 U1619 ( .IN(n2137), .OUT(n558) );
  INVX1 U1620 ( .IN(n2126), .OUT(n569) );
  INVX1 U1621 ( .IN(n2145), .OUT(n552) );
  INVX1 U1622 ( .IN(n2138), .OUT(n557) );
  INVX1 U1623 ( .IN(n2112), .OUT(n583) );
  INVX1 U1624 ( .IN(n2167), .OUT(n531) );
  INVX1 U1625 ( .IN(n2166), .OUT(n532) );
  INVX1 U1626 ( .IN(n2142), .OUT(n553) );
  INVX1 U1627 ( .IN(n2154), .OUT(n544) );
  INVX1 U1628 ( .IN(n2140), .OUT(n555) );
  INVX1 U1629 ( .IN(n2141), .OUT(n554) );
  INVX1 U1630 ( .IN(n2121), .OUT(n574) );
  INVX1 U1631 ( .IN(n2158), .OUT(n540) );
  INVX1 U1632 ( .IN(n2172), .OUT(n526) );
  INVX1 U1633 ( .IN(n2120), .OUT(n575) );
  INVX1 U1634 ( .IN(n2171), .OUT(n527) );
  INVX1 U1635 ( .IN(n2159), .OUT(n539) );
  INVX1 U1636 ( .IN(n2122), .OUT(n573) );
  INVX1 U1637 ( .IN(n2160), .OUT(n538) );
  INVX1 U1638 ( .IN(n2161), .OUT(n537) );
  INVX1 U1639 ( .IN(n2173), .OUT(n525) );
  INVX1 U1640 ( .IN(n2119), .OUT(n576) );
  INVX1 U1641 ( .IN(n2162), .OUT(n536) );
  INVX1 U1642 ( .IN(n2176), .OUT(n522) );
  INVX1 U1643 ( .IN(n2170), .OUT(n528) );
  INVX1 U1644 ( .IN(n2156), .OUT(n542) );
  INVX1 U1645 ( .IN(n2123), .OUT(n572) );
  INVX1 U1646 ( .IN(n2118), .OUT(n577) );
  INVX1 U1647 ( .IN(n2131), .OUT(n564) );
  INVX1 U1648 ( .IN(n2177), .OUT(n521) );
  INVX1 U1649 ( .IN(n2132), .OUT(n563) );
  INVX1 U1650 ( .IN(n2175), .OUT(n523) );
  INVX1 U1651 ( .IN(n2135), .OUT(n560) );
  INVX1 U1652 ( .IN(n2133), .OUT(n562) );
  INVX1 U1653 ( .IN(n2124), .OUT(n571) );
  INVX1 U1654 ( .IN(n2148), .OUT(n550) );
  INVX1 U1655 ( .IN(n2134), .OUT(n561) );
  INVX1 U1656 ( .IN(n2117), .OUT(n578) );
  INVX1 U1657 ( .IN(n2116), .OUT(n579) );
  INVX1 U1658 ( .IN(n2147), .OUT(n551) );
  INVX1 U1659 ( .IN(n2093), .OUT(n596) );
  INVX1 U1660 ( .IN(n2052), .OUT(n702) );
  INVX1 U1661 ( .IN(n2060), .OUT(n700) );
  INVX1 U1662 ( .IN(n2128), .OUT(n567) );
  INVX1 U1663 ( .IN(n2139), .OUT(n556) );
  INVX1 U1664 ( .IN(n2129), .OUT(n566) );
  INVX1 U1665 ( .IN(n2157), .OUT(n541) );
  INVX1 U1666 ( .IN(n2130), .OUT(n565) );
  INVX1 U1667 ( .IN(n2056), .OUT(n701) );
  INVX1 U1668 ( .IN(n2127), .OUT(n568) );
  INVX1 U1669 ( .IN(n2136), .OUT(n559) );
  INVX1 U1670 ( .IN(n2150), .OUT(n548) );
  INVX1 U1671 ( .IN(n2152), .OUT(n546) );
  INVX1 U1672 ( .IN(n2064), .OUT(n699) );
  INVX1 U1673 ( .IN(n2151), .OUT(n547) );
  INVX1 U1674 ( .IN(n2045), .OUT(n2046) );
  INVX1 U1675 ( .IN(n2153), .OUT(n545) );
  INVX1 U1676 ( .IN(n2149), .OUT(n549) );
  INVX1 U1677 ( .IN(n2184), .OUT(n484) );
  INVX1 U1678 ( .IN(n2185), .OUT(n483) );
  INVX1 U1679 ( .IN(n2183), .OUT(n485) );
  NANDX2 U1680 ( .IN1(n1774), .IN2(n1858), .OUT(n2024) );
  INVX1 U1681 ( .IN(n2199), .OUT(n469) );
  INVX1 U1682 ( .IN(n2200), .OUT(n468) );
  INVX1 U1683 ( .IN(n2203), .OUT(n467) );
  BUF4X U1684 ( .IN(n2143), .OUT(n1790) );
  INVX1 U1685 ( .IN(n2197), .OUT(n471) );
  INVX1 U1686 ( .IN(n2196), .OUT(n472) );
  INVX1 U1687 ( .IN(n2195), .OUT(n473) );
  INVX1 U1688 ( .IN(n2198), .OUT(n470) );
  INVX1 U1689 ( .IN(n2194), .OUT(n474) );
  INVX1 U1690 ( .IN(n2193), .OUT(n475) );
  INVX1 U1691 ( .IN(n2190), .OUT(n478) );
  INVX1 U1692 ( .IN(n2192), .OUT(n476) );
  INVX1 U1693 ( .IN(n2186), .OUT(n482) );
  INVX1 U1694 ( .IN(n2187), .OUT(n481) );
  INVX1 U1695 ( .IN(n2191), .OUT(n477) );
  BUF4X U1696 ( .IN(n2179), .OUT(n1793) );
  INVX1 U1697 ( .IN(n2188), .OUT(n480) );
  INVX1 U1698 ( .IN(n2189), .OUT(n479) );
  INVX1 U1699 ( .IN(n2076), .OUT(n614) );
  INVX1 U1700 ( .IN(n2222), .OUT(n414) );
  INVX1 U1701 ( .IN(n2212), .OUT(n424) );
  INVX1 U1702 ( .IN(n2211), .OUT(n425) );
  INVX1 U1703 ( .IN(n2210), .OUT(n426) );
  INVX1 U1704 ( .IN(n2077), .OUT(n613) );
  INVX1 U1705 ( .IN(n2078), .OUT(n612) );
  INVX1 U1706 ( .IN(n2209), .OUT(n427) );
  INVX1 U1707 ( .IN(n2079), .OUT(n611) );
  INVX1 U1708 ( .IN(n2208), .OUT(n428) );
  INVX1 U1709 ( .IN(n2206), .OUT(n430) );
  INVX1 U1710 ( .IN(n2082), .OUT(n610) );
  INVX1 U1711 ( .IN(n2049), .OUT(n2050) );
  INVX1 U1712 ( .IN(n2207), .OUT(n429) );
  INVX1 U1713 ( .IN(n2073), .OUT(n617) );
  INVX1 U1714 ( .IN(n2219), .OUT(n417) );
  INVX1 U1715 ( .IN(n2074), .OUT(n616) );
  NAND2X1 U1716 ( .IN1(n1857), .IN2(n2069), .OUT(n1858) );
  INVX1 U1717 ( .IN(n2220), .OUT(n416) );
  INVX1 U1718 ( .IN(n2218), .OUT(n418) );
  INVX1 U1719 ( .IN(n2214), .OUT(n422) );
  INVX1 U1720 ( .IN(n2221), .OUT(n415) );
  NAND2X1 U1721 ( .IN1(n1979), .IN2(n1978), .OUT(n1980) );
  INVX1 U1722 ( .IN(n2217), .OUT(n419) );
  NAND2X1 U1723 ( .IN1(n1801), .IN2(n1859), .OUT(n1800) );
  INVX1 U1724 ( .IN(n2213), .OUT(n423) );
  INVX1 U1725 ( .IN(n2226), .OUT(n412) );
  INVX1 U1726 ( .IN(n2223), .OUT(n413) );
  INVX1 U1727 ( .IN(n2215), .OUT(n421) );
  INVX1 U1728 ( .IN(n2075), .OUT(n615) );
  INVX1 U1729 ( .IN(n2216), .OUT(n420) );
  NAND2X1 U1730 ( .IN1(n1984), .IN2(n1983), .OUT(n1985) );
  NAND2X1 U1731 ( .IN1(n2204), .IN2(n2181), .OUT(N193) );
  NANDX2 U1732 ( .IN1(n1778), .IN2(n1825), .OUT(n1813) );
  NANDX2 U1733 ( .IN1(n1779), .IN2(n1825), .OUT(n1826) );
  INVX1 U1734 ( .IN(n1860), .OUT(n1857) );
  NANDX2 U1735 ( .IN1(n1777), .IN2(n1825), .OUT(n1822) );
  NANDX2 U1736 ( .IN1(n1775), .IN2(n1825), .OUT(n1816) );
  NANDX2 U1737 ( .IN1(n1776), .IN2(n1825), .OUT(n1819) );
  INVX1 U1738 ( .IN(n1902), .OUT(DEBUG[2]) );
  INVX1 U1739 ( .IN(n1906), .OUT(DEBUG[4]) );
  INVX1 U1740 ( .IN(n1903), .OUT(DEBUG[3]) );
  INVX1 U1741 ( .IN(n1912), .OUT(DOUT[13]) );
  INVX1 U1742 ( .IN(n1925), .OUT(EXC[0]) );
  INVX1 U1743 ( .IN(n1915), .OUT(DOUT[1]) );
  NANDX2 U1744 ( .IN1(n1784), .IN2(Booth_Add_datain1[8]), .OUT(n1877) );
  BUF4X U1745 ( .IN(n2144), .OUT(n1791) );
  INVX1 U1746 ( .IN(n1908), .OUT(DOUT[0]) );
  INVX1 U1747 ( .IN(n1926), .OUT(EXC[1]) );
  INVX1 U1748 ( .IN(n1924), .OUT(DOV) );
  INVX1 U1749 ( .IN(n1894), .OUT(DACK) );
  INVX1 U1750 ( .IN(n1913), .OUT(DOUT[14]) );
  INVX1 U1751 ( .IN(n1927), .OUT(EXC[2]) );
  INVX1 U1752 ( .IN(n1914), .OUT(DOUT[15]) );
  INVX1 U1753 ( .IN(n1922), .OUT(DOUT[8]) );
  INVX1 U1754 ( .IN(n1909), .OUT(DOUT[10]) );
  INVX1 U1755 ( .IN(n1910), .OUT(DOUT[11]) );
  INVX1 U1756 ( .IN(n1921), .OUT(DOUT[7]) );
  INVX1 U1757 ( .IN(AdderCntrl_ExcCheck_Datain[13]), .OUT(n1988) );
  INVX1 U1758 ( .IN(n2053), .OUT(n2054) );
  INVX1 U1759 ( .IN(n1920), .OUT(DOUT[6]) );
  INVX1 U1760 ( .IN(n1923), .OUT(DOUT[9]) );
  INVX1 U1761 ( .IN(n1919), .OUT(DOUT[5]) );
  INVX1 U1762 ( .IN(n1918), .OUT(DOUT[4]) );
  INVX1 U1763 ( .IN(MulCntrl_ExcCheck_Datain[13]), .OUT(n1970) );
  BUF4X U1764 ( .IN(n2178), .OUT(n1792) );
  INVX1 U1765 ( .IN(n1917), .OUT(DOUT[3]) );
  INVX1 U1766 ( .IN(n1911), .OUT(DOUT[12]) );
  INVX1 U1767 ( .IN(n1916), .OUT(DOUT[2]) );
  NAND2X1 U1768 ( .IN1(MulCntrl_ExcCheck_Datain[12]), .IN2(
        MulCntrl_ExcCheck_Datain[11]), .OUT(n1968) );
  NANDX2 U1769 ( .IN1(n1780), .IN2(n1848), .OUT(n1796) );
  INVX1 U1770 ( .IN(n2103), .OUT(n592) );
  NANDX2 U1771 ( .IN1(n1745), .IN2(n1861), .OUT(n1862) );
  INVX1 U1772 ( .IN(n1965), .OUT(n1656) );
  INVX1 U1773 ( .IN(n2020), .OUT(n1587) );
  INVX1 U1774 ( .IN(n2098), .OUT(n594) );
  INVX1 U1775 ( .IN(n1852), .OUT(n1809) );
  INVX1 U1776 ( .IN(n2107), .OUT(n2108) );
  INVX1 U1777 ( .IN(n2057), .OUT(n2058) );
  INVX1 U1778 ( .IN(u_exc_check_N45), .OUT(n2070) );
  INVX1 U1779 ( .IN(n1810), .OUT(n1811) );
  INVX1 U1780 ( .IN(n2099), .OUT(n2101) );
  INVX1 U1781 ( .IN(n2094), .OUT(n2097) );
  INVX1 U1782 ( .IN(n2062), .OUT(n2061) );
  INVX1 U1783 ( .IN(n2036), .OUT(n1964) );
  INVX1 U1784 ( .IN(n2034), .OUT(n2019) );
  INVX1 U1785 ( .IN(n1946), .OUT(n1948) );
  NANDX2 U1786 ( .IN1(multStateMC[0]), .IN2(n1738), .OUT(n1942) );
  NANDX2 U1787 ( .IN1(n462), .IN2(n1744), .OUT(n1946) );
  BUF4X U1788 ( .IN(MulCntrl_Op1[7]), .OUT(n1733) );
  INVX1 U1789 ( .IN(n1895), .OUT(n1901) );
  INVX4 U1790 ( .IN(CS), .OUT(n2029) );
  INVX4 U1791 ( .IN(n1734), .OUT(n1735) );
  INVX4 U1792 ( .IN(RSTn), .OUT(n1795) );
  MUX2X1 U1793 ( .IN1(n1869), .IN2(Add_Op1_wire[0]), .S(n1878), .OUT(
        u_adder_24b_N122) );
  NOR2X1 U1794 ( .IN1(n1869), .IN2(n1878), .OUT(add_x_176_n13) );
  NANDX2 U1795 ( .IN1(n695), .IN2(n694), .OUT(n1807) );
  INVX1 U1796 ( .IN(AdderCntrl_Dataout_valid), .OUT(n1935) );
  NAND2X1 U1797 ( .IN1(n1794), .IN2(n1845), .OUT(n2072) );
  NAND2X1 U1798 ( .IN1(n1794), .IN2(n1966), .OUT(n2107) );
  INVX1 U1799 ( .IN(n2088), .OUT(n600) );
  INVX4 U1800 ( .IN(n1782), .OUT(Booth_ack) );
  INVX8 U1801 ( .IN(n1795), .OUT(n1794) );
  NANDX2 U1802 ( .IN1(n1794), .IN2(n2205), .OUT(n2204) );
  NANDX2 U1803 ( .IN1(n1794), .IN2(n1796), .OUT(n1859) );
  INVX1 U1804 ( .IN(n2091), .OUT(n597) );
  BUF4X U1805 ( .IN(n1886), .OUT(n1784) );
  BUF4X U1806 ( .IN(n1887), .OUT(n1783) );
  INVX4 U1807 ( .IN(n1864), .OUT(n1850) );
  NANDX2 U1808 ( .IN1(n1865), .IN2(n2026), .OUT(n1546) );
  NANDX2 U1809 ( .IN1(n2025), .IN2(n2024), .OUT(n1547) );
  NANDX2 U1810 ( .IN1(n2023), .IN2(n2022), .OUT(n1548) );
  NANDX2 U1811 ( .IN1(n1815), .IN2(n1814), .OUT(n1549) );
  NANDX2 U1812 ( .IN1(n1821), .IN2(n1820), .OUT(n1551) );
  NANDX2 U1813 ( .IN1(n1824), .IN2(n1823), .OUT(n1552) );
  BUF4X U1814 ( .IN(n2201), .OUT(n1788) );
  BUF4X U1815 ( .IN(n1851), .OUT(n1782) );
  BUF4X U1816 ( .IN(n1938), .OUT(n1786) );
  NANDX2 U1817 ( .IN1(n1818), .IN2(n1817), .OUT(n1550) );
  NANDX2 U1818 ( .IN1(n1828), .IN2(n1827), .OUT(n1553) );
  BUF4X U1819 ( .IN(n1941), .OUT(n1785) );
  BUF4X U1820 ( .IN(n2224), .OUT(n1789) );
  INVX4 U1821 ( .IN(n2204), .OUT(n2225) );
  INVX4 U1822 ( .IN(n1859), .OUT(n1855) );
  NANDX2 U1823 ( .IN1(u_exc_check_N45), .IN2(n2004), .OUT(n2005) );
  BUF4X U1824 ( .IN(n2092), .OUT(n1787) );
  NAND2X1 U1825 ( .IN1(u_exc_check_StateMC_0_), .IN2(n1794), .OUT(n2071) );
  NAND2X1 U1826 ( .IN1(n1794), .IN2(n1770), .OUT(n2016) );
  NAND2X1 U1827 ( .IN1(n1748), .IN2(n1794), .OUT(n2035) );
  NAND2X1 U1828 ( .IN1(n1749), .IN2(n1794), .OUT(n2033) );
  NAND2X1 U1829 ( .IN1(n1794), .IN2(Booth_Add_valid), .OUT(n2008) );
  NAND2X1 U1830 ( .IN1(AdderCntrl_ExcCheck_valid), .IN2(n1794), .OUT(n1956) );
  NAND2X1 U1831 ( .IN1(n1794), .IN2(Add_valid), .OUT(n2012) );
  NAND2X1 U1832 ( .IN1(MulCntrl_ExcCheck_valid), .IN2(n1794), .OUT(n1952) );
  INVX1 U1833 ( .IN(MODE[2]), .OUT(n1898) );
  NAND2X1 U1834 ( .IN1(n1794), .IN2(n1936), .OUT(n1937) );
  INVX4 U1835 ( .IN(n1813), .OUT(u_booth_N53) );
  INVX4 U1836 ( .IN(n1816), .OUT(u_booth_N52) );
  INVX4 U1837 ( .IN(n1826), .OUT(u_booth_N49) );
  INVX4 U1838 ( .IN(n1819), .OUT(u_booth_N51) );
  INVX4 U1839 ( .IN(n1822), .OUT(u_booth_N50) );
  INVX4 U1840 ( .IN(n2072), .OUT(n2080) );
  NANDX2 U1841 ( .IN1(n1864), .IN2(n1863), .OUT(n2081) );
  NAND2X1 U1842 ( .IN1(n1794), .IN2(u_booth_BStateMC_1_), .OUT(n1864) );
  NAND2X1 U1843 ( .IN1(n1794), .IN2(n1939), .OUT(n1940) );
  NAND2X1 U1844 ( .IN1(n587), .IN2(CS), .OUT(n1907) );
  NANDX2 U1845 ( .IN1(n1868), .IN2(n1861), .OUT(n1812) );
  INVX4 U1846 ( .IN(n1804), .OUT(n1856) );
  INVX4 U1847 ( .IN(n2043), .OUT(n2065) );
  INVX4 U1848 ( .IN(n2021), .OUT(n1868) );
  NANDX2 U1849 ( .IN1(n1798), .IN2(n1861), .OUT(n1804) );
  NANDX2 U1850 ( .IN1(n2040), .IN2(n2039), .OUT(n2044) );
  INVX4 U1851 ( .IN(n1862), .OUT(n2040) );
  NAND2X1 U1852 ( .IN1(n1794), .IN2(n1830), .OUT(n1797) );
  INVX4 U1853 ( .IN(n2105), .OUT(n2003) );
  NANDX2 U1854 ( .IN1(n1993), .IN2(n1998), .OUT(n2105) );
  INVX4 U1855 ( .IN(n1869), .OUT(Add_Op1_wire[0]) );
  INVX4 U1856 ( .IN(n1879), .OUT(Add_Op2_wire[1]) );
  INVX4 U1857 ( .IN(n1870), .OUT(Add_Op1_wire[1]) );
  INVX4 U1858 ( .IN(n1880), .OUT(Add_Op2_wire[2]) );
  INVX4 U1859 ( .IN(n1871), .OUT(Add_Op1_wire[2]) );
  INVX4 U1860 ( .IN(n1881), .OUT(Add_Op2_wire[3]) );
  INVX4 U1861 ( .IN(n1872), .OUT(Add_Op1_wire[3]) );
  INVX4 U1862 ( .IN(n1882), .OUT(Add_Op2_wire[4]) );
  INVX4 U1863 ( .IN(n1873), .OUT(Add_Op1_wire[4]) );
  INVX4 U1864 ( .IN(n1883), .OUT(Add_Op2_wire[5]) );
  INVX4 U1865 ( .IN(n1874), .OUT(Add_Op1_wire[5]) );
  INVX4 U1866 ( .IN(n1884), .OUT(Add_Op2_wire[6]) );
  INVX4 U1867 ( .IN(n1875), .OUT(Add_Op1_wire[6]) );
  INVX4 U1868 ( .IN(n1885), .OUT(Add_Op2_wire[7]) );
  INVX4 U1869 ( .IN(n1876), .OUT(Add_Op1_wire[7]) );
  INVX4 U1870 ( .IN(n1888), .OUT(Add_Op2_wire[8]) );
  INVX4 U1871 ( .IN(n1877), .OUT(Add_Op1_wire[8]) );
  NAND2X1 U1872 ( .IN1(n1773), .IN2(n1858), .OUT(n2022) );
  INVX4 U1873 ( .IN(n2044), .OUT(n2066) );
  INVX4 U1874 ( .IN(n1942), .OUT(n2182) );
  NAND2X1 U1875 ( .IN1(n2021), .IN2(n1745), .OUT(n1798) );
  TIEHI U1876 ( .OUT(n408) );
  NAND2X1 U1877 ( .IN1(n1810), .IN2(n1861), .OUT(n1808) );
  NAND2X1 U1878 ( .IN1(u_booth_count_reg_2_), .IN2(n1855), .OUT(n1802) );
  NAND2X1 U1879 ( .IN1(u_booth_count_reg_2_), .IN2(n1801), .OUT(n1805) );
  INVX4 U1880 ( .IN(n2038), .OUT(u_adder_24b_N52) );
  INVX4 U1881 ( .IN(n2181), .OUT(n2202) );
  NOR2X1 U1882 ( .IN1(u_booth_BStateMC_1_), .IN2(n1781), .OUT(n1853) );
  AOI22 U1883 ( .IN1(n1830), .IN2(n2006), .IN3(Booth_valid), .IN4(n1853), 
        .OUT(n1848) );
  INVX4 U1884 ( .IN(n1797), .OUT(n1861) );
  MUX2X1 U1885 ( .IN1(n1855), .IN2(n1856), .S(n694), .OUT(n1554) );
  NOR2X1 U1886 ( .IN1(n694), .IN2(n695), .OUT(n1801) );
  OAI21 U1887 ( .IN1(n695), .IN2(n1859), .IN3(n1804), .OUT(n1799) );
  NAND3X1 U1888 ( .IN1(n1807), .IN2(n1800), .IN3(n1799), .OUT(n1079) );
  OAI21 U1889 ( .IN1(n1801), .IN2(u_booth_count_reg_2_), .IN3(n1805), .OUT(
        n1803) );
  OAI21 U1890 ( .IN1(n1804), .IN2(n1803), .IN3(n1802), .OUT(n1555) );
  MUX2X1 U1891 ( .IN1(n1767), .IN2(u_booth_count_reg_3_), .S(n1805), .OUT(
        n1806) );
  AOI22 U1892 ( .IN1(n1856), .IN2(n1806), .IN3(u_booth_count_reg_3_), .IN4(
        n1855), .OUT(n1092) );
  NOR2X1 U1893 ( .IN1(n732), .IN2(n1864), .OUT(n1852) );
  OAI21 U1894 ( .IN1(u_booth_count_reg_2_), .IN2(n1807), .IN3(
        u_booth_count_reg_3_), .OUT(n1810) );
  NAND3X1 U1895 ( .IN1(n1809), .IN2(n1808), .IN3(n2072), .OUT(n1556) );
  NANDX2 U1896 ( .IN1(n1830), .IN2(n1811), .OUT(n1851) );
  AOI21 U1897 ( .IN1(Booth_ack), .IN2(n1794), .IN3(n1852), .OUT(n1088) );
  NANDX2 U1898 ( .IN1(n2006), .IN2(n1861), .OUT(n2069) );
  AOI22 U1899 ( .IN1(n1778), .IN2(n1860), .IN3(Add_dataout[5]), .IN4(n1866), 
        .OUT(n1815) );
  INVX4 U1900 ( .IN(n1812), .OUT(n1867) );
  INVX4 U1901 ( .IN(n2069), .OUT(n1825) );
  AOI21 U1902 ( .IN1(n1867), .IN2(n1773), .IN3(u_booth_N53), .OUT(n1814) );
  AOI22 U1903 ( .IN1(n1860), .IN2(n1775), .IN3(Add_dataout[4]), .IN4(n1866), 
        .OUT(n1818) );
  AOI21 U1904 ( .IN1(n1867), .IN2(n1778), .IN3(u_booth_N52), .OUT(n1817) );
  AOI22 U1905 ( .IN1(n1860), .IN2(n1776), .IN3(Add_dataout[3]), .IN4(n1866), 
        .OUT(n1821) );
  AOI21 U1906 ( .IN1(n1867), .IN2(n1775), .IN3(u_booth_N51), .OUT(n1820) );
  AOI22 U1907 ( .IN1(n1860), .IN2(n1777), .IN3(Add_dataout[2]), .IN4(n1866), 
        .OUT(n1824) );
  AOI21 U1908 ( .IN1(n1867), .IN2(n1776), .IN3(u_booth_N50), .OUT(n1823) );
  AOI22 U1909 ( .IN1(n1779), .IN2(n1860), .IN3(Add_dataout[1]), .IN4(n1866), 
        .OUT(n1828) );
  AOI21 U1910 ( .IN1(n1867), .IN2(n1777), .IN3(u_booth_N49), .OUT(n1827) );
  AOI22 U1911 ( .IN1(n1867), .IN2(n1779), .IN3(n1866), .IN4(Add_dataout[0]), 
        .OUT(n1829) );
  OAI21 U1912 ( .IN1(n721), .IN2(n1859), .IN3(n1829), .OUT(n1544) );
  AOI22 U1913 ( .IN1(n1846), .IN2(n1768), .IN3(Booth_datain2[7]), .IN4(n1845), 
        .OUT(n1831) );
  OAI21 U1914 ( .IN1(n1848), .IN2(n720), .IN3(n1831), .OUT(n1832) );
  AOI22 U1915 ( .IN1(n1850), .IN2(n1759), .IN3(n1794), .IN4(n1832), .OUT(n1022) );
  AOI22 U1916 ( .IN1(n1846), .IN2(n1759), .IN3(Booth_datain2[6]), .IN4(n1845), 
        .OUT(n1833) );
  OAI21 U1917 ( .IN1(n1848), .IN2(n719), .IN3(n1833), .OUT(n1834) );
  AOI22 U1918 ( .IN1(n1850), .IN2(n1760), .IN3(n1794), .IN4(n1834), .OUT(n1028) );
  AOI22 U1919 ( .IN1(n1846), .IN2(n1760), .IN3(Booth_datain2[5]), .IN4(n1845), 
        .OUT(n1835) );
  OAI21 U1920 ( .IN1(n1848), .IN2(n718), .IN3(n1835), .OUT(n1836) );
  AOI22 U1921 ( .IN1(n1850), .IN2(n1761), .IN3(n1794), .IN4(n1836), .OUT(n1031) );
  AOI22 U1922 ( .IN1(n1846), .IN2(n1761), .IN3(Booth_datain2[4]), .IN4(n1845), 
        .OUT(n1837) );
  OAI21 U1923 ( .IN1(n1848), .IN2(n717), .IN3(n1837), .OUT(n1838) );
  AOI22 U1924 ( .IN1(n1850), .IN2(n1762), .IN3(n1794), .IN4(n1838), .OUT(n1034) );
  AOI22 U1925 ( .IN1(n1846), .IN2(n1762), .IN3(Booth_datain2[3]), .IN4(n1845), 
        .OUT(n1839) );
  OAI21 U1926 ( .IN1(n1848), .IN2(n716), .IN3(n1839), .OUT(n1840) );
  AOI22 U1927 ( .IN1(n1850), .IN2(n1763), .IN3(n1794), .IN4(n1840), .OUT(n1037) );
  AOI22 U1928 ( .IN1(n1846), .IN2(n1763), .IN3(Booth_datain2[2]), .IN4(n1845), 
        .OUT(n1841) );
  OAI21 U1929 ( .IN1(n1848), .IN2(n715), .IN3(n1841), .OUT(n1842) );
  AOI22 U1930 ( .IN1(n1850), .IN2(n1764), .IN3(n1794), .IN4(n1842), .OUT(n1040) );
  AOI22 U1931 ( .IN1(n1846), .IN2(n1764), .IN3(Booth_datain2[1]), .IN4(n1845), 
        .OUT(n1843) );
  OAI21 U1932 ( .IN1(n1848), .IN2(n714), .IN3(n1843), .OUT(n1844) );
  AOI22 U1933 ( .IN1(n1850), .IN2(n1765), .IN3(n1794), .IN4(n1844), .OUT(n1043) );
  AOI22 U1934 ( .IN1(n1846), .IN2(n1765), .IN3(Booth_datain2[0]), .IN4(n1845), 
        .OUT(n1847) );
  OAI21 U1935 ( .IN1(n1848), .IN2(n713), .IN3(n1847), .OUT(n1849) );
  AOI22 U1936 ( .IN1(n1850), .IN2(n1736), .IN3(n1794), .IN4(n1849), .OUT(n1135) );
  NOR2X1 U1937 ( .IN1(n713), .IN2(n1782), .OUT(Booth_dataout[0]) );
  NOR2X1 U1938 ( .IN1(n714), .IN2(n1782), .OUT(Booth_dataout[1]) );
  NOR2X1 U1939 ( .IN1(n715), .IN2(n1782), .OUT(Booth_dataout[2]) );
  NOR2X1 U1940 ( .IN1(n716), .IN2(n1851), .OUT(Booth_dataout[3]) );
  NOR2X1 U1941 ( .IN1(n717), .IN2(n1851), .OUT(Booth_dataout[4]) );
  NOR2X1 U1942 ( .IN1(n718), .IN2(n1851), .OUT(Booth_dataout[5]) );
  NOR2X1 U1943 ( .IN1(n719), .IN2(n1851), .OUT(Booth_dataout[6]) );
  NOR2X1 U1944 ( .IN1(n720), .IN2(n1851), .OUT(Booth_dataout[7]) );
  NOR2X1 U1945 ( .IN1(n721), .IN2(n1851), .OUT(Booth_dataout[8]) );
  NOR2X1 U1946 ( .IN1(n722), .IN2(n1851), .OUT(Booth_dataout[9]) );
  NOR2X1 U1947 ( .IN1(n723), .IN2(n1851), .OUT(Booth_dataout[10]) );
  NOR2X1 U1948 ( .IN1(n724), .IN2(n1851), .OUT(Booth_dataout[11]) );
  NOR2X1 U1949 ( .IN1(n725), .IN2(n1851), .OUT(Booth_dataout[12]) );
  NOR2X1 U1950 ( .IN1(n726), .IN2(n1851), .OUT(Booth_dataout[13]) );
  NOR2X1 U1951 ( .IN1(n727), .IN2(n1782), .OUT(Booth_dataout[14]) );
  NOR2X1 U1952 ( .IN1(n728), .IN2(n1782), .OUT(Booth_dataout[15]) );
  AOI21 U1953 ( .IN1(n1853), .IN2(n1794), .IN3(n1852), .OUT(n1854) );
  OAI21 U1954 ( .IN1(n1854), .IN2(n1758), .IN3(n2069), .OUT(n1653) );
  AOI22 U1955 ( .IN1(n1856), .IN2(n1736), .IN3(u_booth_Q1_reg), .IN4(n1855), 
        .OUT(n1077) );
  AOI22 U1956 ( .IN1(n1867), .IN2(u_booth_A_reg_8_), .IN3(n1866), .IN4(
        Add_dataout[8]), .OUT(n1865) );
  OAI21 U1957 ( .IN1(n1859), .IN2(n1771), .IN3(n1865), .OUT(n1545) );
  NOR2X1 U1958 ( .IN1(n1756), .IN2(n2069), .OUT(n706) );
  AOI21 U1959 ( .IN1(u_booth_A_reg_7_), .IN2(n1860), .IN3(n706), .OUT(n2026)
         );
  OAI21 U1960 ( .IN1(Booth_valid), .IN2(n1781), .IN3(n1794), .OUT(n1863) );
  NOR2X1 U1961 ( .IN1(n728), .IN2(n2069), .OUT(u_booth_N55) );
  NOR2X1 U1962 ( .IN1(n727), .IN2(n2069), .OUT(u_booth_N54) );
  NOR2X1 U1963 ( .IN1(AddSelect), .IN2(n802), .OUT(n1887) );
  NOR2X1 U1964 ( .IN1(n802), .IN2(n1783), .OUT(n1886) );
  AOI22 U1965 ( .IN1(n1783), .IN2(Add_Op1[0]), .IN3(n1784), .IN4(
        Booth_Add_datain1[0]), .OUT(n1869) );
  AOI22 U1966 ( .IN1(n1783), .IN2(Add_Op1[1]), .IN3(n1784), .IN4(
        Booth_Add_datain1[1]), .OUT(n1870) );
  AOI22 U1967 ( .IN1(n1783), .IN2(Add_Op1[2]), .IN3(n1784), .IN4(
        Booth_Add_datain1[2]), .OUT(n1871) );
  AOI22 U1968 ( .IN1(n1783), .IN2(Add_Op1[3]), .IN3(n1784), .IN4(
        Booth_Add_datain1[3]), .OUT(n1872) );
  AOI22 U1969 ( .IN1(n1783), .IN2(Add_Op1[4]), .IN3(n1784), .IN4(
        Booth_Add_datain1[4]), .OUT(n1873) );
  AOI22 U1970 ( .IN1(n1783), .IN2(Add_Op1[5]), .IN3(n1784), .IN4(
        Booth_Add_datain1[5]), .OUT(n1874) );
  AOI22 U1971 ( .IN1(n1783), .IN2(Add_Op1[6]), .IN3(n1784), .IN4(
        Booth_Add_datain1[6]), .OUT(n1875) );
  AOI22 U1972 ( .IN1(n1783), .IN2(Add_Op1[7]), .IN3(n1784), .IN4(
        Booth_Add_datain1[7]), .OUT(n1876) );
  AOI22 U1973 ( .IN1(n1783), .IN2(Add_Op2[0]), .IN3(n1784), .IN4(
        Booth_Add_datain2[0]), .OUT(n1878) );
  AOI22 U1974 ( .IN1(n1783), .IN2(Add_Op2[1]), .IN3(n1784), .IN4(
        Booth_Add_datain2[1]), .OUT(n1879) );
  AOI22 U1975 ( .IN1(n1783), .IN2(Add_Op2[2]), .IN3(n1784), .IN4(
        Booth_Add_datain2[2]), .OUT(n1880) );
  AOI22 U1976 ( .IN1(n1783), .IN2(Add_Op2[3]), .IN3(n1784), .IN4(
        Booth_Add_datain2[3]), .OUT(n1881) );
  AOI22 U1977 ( .IN1(n1783), .IN2(Add_Op2[4]), .IN3(n1784), .IN4(
        Booth_Add_datain2[4]), .OUT(n1882) );
  AOI22 U1978 ( .IN1(n1783), .IN2(Add_Op2[5]), .IN3(n1784), .IN4(
        Booth_Add_datain2[5]), .OUT(n1883) );
  AOI22 U1979 ( .IN1(n1783), .IN2(Add_Op2[6]), .IN3(n1784), .IN4(
        Booth_Add_datain2[6]), .OUT(n1884) );
  AOI22 U1980 ( .IN1(n1783), .IN2(Add_Op2[7]), .IN3(n1784), .IN4(
        Booth_Add_datain2[7]), .OUT(n1885) );
  AOI22 U1981 ( .IN1(n1783), .IN2(Add_Op2[8]), .IN3(n1784), .IN4(
        Booth_Add_datain2[8]), .OUT(n1888) );
  NAND3X1 U1982 ( .IN1(getdataStat_reg[0]), .IN2(n463), .IN3(ABUSY), .OUT(
        n1889) );
  NOR2X1 U1983 ( .IN1(n1889), .IN2(n1741), .OUT(AdderCntrl_valid) );
  NOR2X1 U1984 ( .IN1(ABUSY), .IN2(OPT), .OUT(n1890) );
  NAND3X1 U1985 ( .IN1(CS), .IN2(DIV), .IN3(n1890), .OUT(n1891) );
  NOR2X1 U1986 ( .IN1(getdataStat_reg[0]), .IN2(n1891), .OUT(n2146) );
  NOR2X1 U1987 ( .IN1(MBUSY), .IN2(getdataStat_reg[1]), .OUT(n1892) );
  NAND3X1 U1988 ( .IN1(DIV), .IN2(OPT), .IN3(n1892), .OUT(n1893) );
  NOR2X1 U1989 ( .IN1(n2029), .IN2(n1893), .OUT(n2111) );
  NOR2X1 U1990 ( .IN1(n2146), .IN2(n2111), .OUT(n1894) );
  NOR2X1 U1991 ( .IN1(MODE[1]), .IN2(MODE[0]), .OUT(n1895) );
  AOI22 U1992 ( .IN1(MODE[2]), .IN2(multStateMC[0]), .IN3(n1744), .IN4(n1898), 
        .OUT(n1897) );
  NOR2X1 U1993 ( .IN1(n1895), .IN2(MODE[2]), .OUT(n1905) );
  NOR2X1 U1994 ( .IN1(n1895), .IN2(n1898), .OUT(n1904) );
  AOI22 U1995 ( .IN1(n1905), .IN2(AdderCntrl_Debug[0]), .IN3(n1904), .IN4(
        MulCntrl_Debug[0]), .OUT(n1896) );
  OAI21 U1996 ( .IN1(n1901), .IN2(n1897), .IN3(n1896), .OUT(DEBUG[0]) );
  AOI22 U1997 ( .IN1(MODE[2]), .IN2(multStateMC[1]), .IN3(n1741), .IN4(n1898), 
        .OUT(n1900) );
  AOI22 U1998 ( .IN1(n1905), .IN2(AdderCntrl_Debug[1]), .IN3(n1904), .IN4(
        MulCntrl_Debug[1]), .OUT(n1899) );
  OAI21 U1999 ( .IN1(n1901), .IN2(n1900), .IN3(n1899), .OUT(DEBUG[1]) );
  AOI22 U2000 ( .IN1(n1905), .IN2(AdderCntrl_Debug[2]), .IN3(n1904), .IN4(
        MulCntrl_Debug[2]), .OUT(n1902) );
  AOI22 U2001 ( .IN1(n1905), .IN2(AdderCntrl_Debug[3]), .IN3(n1904), .IN4(
        MulCntrl_Debug[3]), .OUT(n1903) );
  AOI22 U2002 ( .IN1(n1905), .IN2(AdderCntrl_Debug[4]), .IN3(n1904), .IN4(
        MulCntrl_Debug[4]), .OUT(n1906) );
  NOR2X1 U2003 ( .IN1(n584), .IN2(n1907), .OUT(n1941) );
  NOR2X1 U2004 ( .IN1(n587), .IN2(n2029), .OUT(n1938) );
  AOI22 U2005 ( .IN1(n1785), .IN2(MultResult_reg[0]), .IN3(AdderResult_reg[0]), 
        .IN4(n1786), .OUT(n1908) );
  AOI22 U2006 ( .IN1(n1785), .IN2(MultResult_reg[10]), .IN3(
        AdderResult_reg[10]), .IN4(n1786), .OUT(n1909) );
  AOI22 U2007 ( .IN1(n1785), .IN2(MultResult_reg[11]), .IN3(
        AdderResult_reg[11]), .IN4(n1786), .OUT(n1910) );
  AOI22 U2008 ( .IN1(n1785), .IN2(MultResult_reg[12]), .IN3(
        AdderResult_reg[12]), .IN4(n1786), .OUT(n1911) );
  AOI22 U2009 ( .IN1(n1785), .IN2(MultResult_reg[13]), .IN3(
        AdderResult_reg[13]), .IN4(n1786), .OUT(n1912) );
  AOI22 U2010 ( .IN1(n1785), .IN2(MultResult_reg[14]), .IN3(
        AdderResult_reg[14]), .IN4(n1786), .OUT(n1913) );
  AOI22 U2011 ( .IN1(n1785), .IN2(MultResult_reg[15]), .IN3(
        AdderResult_reg[15]), .IN4(n1786), .OUT(n1914) );
  AOI22 U2012 ( .IN1(n1785), .IN2(MultResult_reg[1]), .IN3(AdderResult_reg[1]), 
        .IN4(n1786), .OUT(n1915) );
  AOI22 U2013 ( .IN1(n1785), .IN2(MultResult_reg[2]), .IN3(AdderResult_reg[2]), 
        .IN4(n1786), .OUT(n1916) );
  AOI22 U2014 ( .IN1(n1785), .IN2(MultResult_reg[3]), .IN3(AdderResult_reg[3]), 
        .IN4(n1786), .OUT(n1917) );
  AOI22 U2015 ( .IN1(n1785), .IN2(MultResult_reg[4]), .IN3(AdderResult_reg[4]), 
        .IN4(n1786), .OUT(n1918) );
  AOI22 U2016 ( .IN1(n1785), .IN2(MultResult_reg[5]), .IN3(AdderResult_reg[5]), 
        .IN4(n1786), .OUT(n1919) );
  AOI22 U2017 ( .IN1(n1785), .IN2(MultResult_reg[6]), .IN3(AdderResult_reg[6]), 
        .IN4(n1786), .OUT(n1920) );
  AOI22 U2018 ( .IN1(n1785), .IN2(MultResult_reg[7]), .IN3(AdderResult_reg[7]), 
        .IN4(n1786), .OUT(n1921) );
  AOI22 U2019 ( .IN1(n1785), .IN2(MultResult_reg[8]), .IN3(AdderResult_reg[8]), 
        .IN4(n1786), .OUT(n1922) );
  AOI22 U2020 ( .IN1(n1785), .IN2(MultResult_reg[9]), .IN3(AdderResult_reg[9]), 
        .IN4(n1786), .OUT(n1923) );
  NOR2X1 U2021 ( .IN1(n1785), .IN2(n1786), .OUT(n1924) );
  AOI22 U2022 ( .IN1(n1785), .IN2(MultExc_reg[0]), .IN3(AddExc_reg[0]), .IN4(
        n1786), .OUT(n1925) );
  AOI22 U2023 ( .IN1(n1785), .IN2(MultExc_reg[1]), .IN3(AddExc_reg[1]), .IN4(
        n1786), .OUT(n1926) );
  AOI22 U2024 ( .IN1(n1785), .IN2(MultExc_reg[2]), .IN3(AddExc_reg[2]), .IN4(
        n1786), .OUT(n1927) );
  NAND3X1 U2025 ( .IN1(getdataStat_reg[1]), .IN2(MBUSY), .IN3(n1746), .OUT(
        n1928) );
  NOR2X1 U2026 ( .IN1(multStateMC[1]), .IN2(n1928), .OUT(MulCntrl_valid) );
  NAND3X1 U2027 ( .IN1(n463), .IN2(n587), .IN3(n1741), .OUT(n1931) );
  OAI21 U2028 ( .IN1(getdataStat_reg[0]), .IN2(n2146), .IN3(n1931), .OUT(n1929) );
  NOR2X1 U2029 ( .IN1(n1795), .IN2(n1929), .OUT(N149) );
  NAND3X1 U2030 ( .IN1(multStateMC[1]), .IN2(n584), .IN3(n1746), .OUT(n1933)
         );
  OAI21 U2031 ( .IN1(getdataStat_reg[1]), .IN2(n2111), .IN3(n1933), .OUT(n1930) );
  NOR2X1 U2032 ( .IN1(n1795), .IN2(n1930), .OUT(N150) );
  OAI21 U2033 ( .IN1(ABUSY), .IN2(n2146), .IN3(n1931), .OUT(n1932) );
  AOI21 U2034 ( .IN1(n1946), .IN2(n1932), .IN3(n1795), .OUT(N151) );
  OAI21 U2035 ( .IN1(MBUSY), .IN2(n2111), .IN3(n1933), .OUT(n1934) );
  AOI21 U2036 ( .IN1(n1942), .IN2(n1934), .IN3(n1795), .OUT(N152) );
  NAND2X1 U2037 ( .IN1(CS), .IN2(n1935), .OUT(n1947) );
  OAI21 U2038 ( .IN1(n1947), .IN2(n1946), .IN3(n587), .OUT(n1936) );
  AOI21 U2039 ( .IN1(DOA), .IN2(n1786), .IN3(n1937), .OUT(N191) );
  NAND2X1 U2040 ( .IN1(CS), .IN2(MulCntrl_Dataout_valid), .OUT(n2030) );
  OAI21 U2041 ( .IN1(n2030), .IN2(n1942), .IN3(n584), .OUT(n1939) );
  AOI21 U2042 ( .IN1(n1785), .IN2(DOA), .IN3(n1940), .OUT(N192) );
  NOR2X1 U2043 ( .IN1(AdderCntrl_Dataout_valid), .IN2(n1946), .OUT(n2205) );
  NAND3X1 U2044 ( .IN1(n1794), .IN2(n2182), .IN3(MulCntrl_Dataout_valid), 
        .OUT(n2181) );
  NAND3X1 U2045 ( .IN1(n806), .IN2(u_Adder_interconnect_stateMC_1_), .IN3(
        Booth_Add_valid), .OUT(n2034) );
  NAND3X1 U2046 ( .IN1(Add_valid), .IN2(n1739), .IN3(n1754), .OUT(n2094) );
  NAND2X1 U2047 ( .IN1(AddSelect), .IN2(n2094), .OUT(n1943) );
  AOI21 U2048 ( .IN1(n2034), .IN2(n1943), .IN3(n1795), .OUT(n1723) );
  AOI21 U2049 ( .IN1(n587), .IN2(n463), .IN3(n1795), .OUT(n1944) );
  NAND2X1 U2050 ( .IN1(n1741), .IN2(n1944), .OUT(n1945) );
  OAI21 U2051 ( .IN1(n2029), .IN2(n2204), .IN3(n1945), .OUT(n1692) );
  AOI21 U2052 ( .IN1(n1948), .IN2(n1947), .IN3(AdderCntrl_valid), .OUT(n1949)
         );
  OAI21 U2053 ( .IN1(n463), .IN2(n462), .IN3(n1949), .OUT(n1950) );
  NAND2X1 U2054 ( .IN1(n1794), .IN2(n1950), .OUT(n1302) );
  NOR2X1 U2055 ( .IN1(u_ExcChecker_interconnect_stateMC_0_), .IN2(
        u_ExcChecker_interconnect_stateMC_1_), .OUT(n1963) );
  NAND2X1 U2056 ( .IN1(AdderCntrl_ExcCheck_valid), .IN2(n1752), .OUT(n1951) );
  AOI22 U2057 ( .IN1(u_ExcChecker_interconnect_stateMC_1_), .IN2(n1748), .IN3(
        n1963), .IN4(n1951), .OUT(n1953) );
  NAND3X1 U2058 ( .IN1(n1794), .IN2(u_ExcChecker_interconnect_stateMC_0_), 
        .IN3(u_ExcChecker_interconnect_stateMC_1_), .OUT(n1955) );
  OAI21 U2059 ( .IN1(n1953), .IN2(n1952), .IN3(n1955), .OUT(n1661) );
  NAND2X1 U2060 ( .IN1(MulCntrl_ExcCheck_valid), .IN2(
        u_ExcChecker_interconnect_priority_reg), .OUT(n1954) );
  AOI22 U2061 ( .IN1(u_ExcChecker_interconnect_stateMC_0_), .IN2(n1748), .IN3(
        n1963), .IN4(n1954), .OUT(n1957) );
  OAI21 U2062 ( .IN1(n1957), .IN2(n1956), .IN3(n1955), .OUT(n1660) );
  INVX1 U2063 ( .IN(MulCntrl_ExcCheck_valid), .OUT(n1958) );
  AOI22 U2064 ( .IN1(u_ExcChecker_interconnect_priority_reg), .IN2(n1958), 
        .IN3(AdderCntrl_ExcCheck_valid), .IN4(n1752), .OUT(n1960) );
  OAI21 U2065 ( .IN1(u_ExcChecker_interconnect_priority_reg), .IN2(n1963), 
        .IN3(n1794), .OUT(n1959) );
  AOI21 U2066 ( .IN1(n1963), .IN2(n1960), .IN3(n1959), .OUT(n1659) );
  NAND3X1 U2067 ( .IN1(u_ExcChecker_interconnect_stateMC_1_), .IN2(
        MulCntrl_ExcCheck_valid), .IN3(n1753), .OUT(n2036) );
  NAND3X1 U2068 ( .IN1(u_ExcChecker_interconnect_stateMC_0_), .IN2(
        AdderCntrl_ExcCheck_valid), .IN3(n1755), .OUT(n2099) );
  NAND2X1 U2069 ( .IN1(ExcSelect), .IN2(n2099), .OUT(n1961) );
  AOI21 U2070 ( .IN1(n2036), .IN2(n1961), .IN3(n1795), .OUT(n1658) );
  AOI21 U2071 ( .IN1(ExcCheck_valid), .IN2(n1772), .IN3(u_exc_check_StateMC_0_), .OUT(n1962) );
  NOR2X1 U2072 ( .IN1(n1962), .IN2(n1795), .OUT(n1657) );
  NAND3X1 U2073 ( .IN1(n654), .IN2(ExcCheck_valid), .IN3(n1766), .OUT(n1966)
         );
  NOR2X1 U2074 ( .IN1(n1795), .IN2(n1966), .OUT(u_exc_check_N45) );
  NOR2X1 U2075 ( .IN1(n1963), .IN2(n1795), .OUT(n2102) );
  NOR2X1 U2076 ( .IN1(n1795), .IN2(n1748), .OUT(n2100) );
  AOI22 U2077 ( .IN1(n2102), .IN2(MulCntrl_Exc_Ack), .IN3(n1964), .IN4(n2100), 
        .OUT(n1965) );
  NAND3X1 U2078 ( .IN1(MulCntrl_ExcCheck_Datain[10]), .IN2(
        MulCntrl_ExcCheck_Datain[7]), .IN3(ExcSelect), .OUT(n1967) );
  NOR2X1 U2079 ( .IN1(n1968), .IN2(n1967), .OUT(n1977) );
  NAND3X1 U2080 ( .IN1(MulCntrl_ExcCheck_Datain[14]), .IN2(
        MulCntrl_ExcCheck_Datain[8]), .IN3(MulCntrl_ExcCheck_Datain[9]), .OUT(
        n1969) );
  NOR2X1 U2081 ( .IN1(n1970), .IN2(n1969), .OUT(n1976) );
  NOR2X1 U2082 ( .IN1(AdderCntrl_ExcCheck_Datain[13]), .IN2(
        AdderCntrl_ExcCheck_Datain[10]), .OUT(n1971) );
  NAND3X1 U2083 ( .IN1(n1971), .IN2(AdderCntrl_ExcCheck_Datain[8]), .IN3(
        AdderCntrl_ExcCheck_Datain[9]), .OUT(n1972) );
  NOR2X1 U2084 ( .IN1(ExcSelect), .IN2(n1972), .OUT(n1975) );
  NAND3X1 U2085 ( .IN1(AdderCntrl_ExcCheck_Datain[11]), .IN2(
        AdderCntrl_ExcCheck_Datain[12]), .IN3(AdderCntrl_ExcCheck_Datain[14]), 
        .OUT(n1973) );
  NOR2X1 U2086 ( .IN1(AdderCntrl_ExcCheck_Datain[7]), .IN2(n1973), .OUT(n1974)
         );
  AOI22 U2087 ( .IN1(n1977), .IN2(n1976), .IN3(n1975), .IN4(n1974), .OUT(n2106) );
  NOR2X1 U2088 ( .IN1(AdderCntrl_ExcCheck_Datain[3]), .IN2(
        AdderCntrl_ExcCheck_Datain[4]), .OUT(n1979) );
  NOR2X1 U2089 ( .IN1(AdderCntrl_ExcCheck_Datain[2]), .IN2(
        AdderCntrl_ExcCheck_Datain[0]), .OUT(n1978) );
  NOR2X1 U2090 ( .IN1(AdderCntrl_ExcCheck_Datain[1]), .IN2(n1980), .OUT(n1982)
         );
  NOR2X1 U2091 ( .IN1(AdderCntrl_ExcCheck_Datain[5]), .IN2(
        AdderCntrl_ExcCheck_Datain[6]), .OUT(n1981) );
  NAND3X1 U2092 ( .IN1(n1982), .IN2(n1981), .IN3(n1747), .OUT(n1993) );
  NOR2X1 U2093 ( .IN1(MulCntrl_ExcCheck_Datain[3]), .IN2(
        MulCntrl_ExcCheck_Datain[4]), .OUT(n1984) );
  NOR2X1 U2094 ( .IN1(MulCntrl_ExcCheck_Datain[2]), .IN2(
        MulCntrl_ExcCheck_Datain[0]), .OUT(n1983) );
  NOR2X1 U2095 ( .IN1(MulCntrl_ExcCheck_Datain[1]), .IN2(n1985), .OUT(n1987)
         );
  NOR2X1 U2096 ( .IN1(MulCntrl_ExcCheck_Datain[5]), .IN2(
        MulCntrl_ExcCheck_Datain[6]), .OUT(n1986) );
  NAND3X1 U2097 ( .IN1(n1987), .IN2(n1986), .IN3(ExcSelect), .OUT(n1998) );
  NOR2X1 U2098 ( .IN1(AdderCntrl_ExcCheck_Datain[14]), .IN2(
        AdderCntrl_ExcCheck_Datain[9]), .OUT(n2002) );
  NOR2X1 U2099 ( .IN1(AdderCntrl_ExcCheck_Datain[12]), .IN2(n1988), .OUT(n1991) );
  NOR2X1 U2100 ( .IN1(AdderCntrl_ExcCheck_Datain[11]), .IN2(n1731), .OUT(n1990) );
  NOR2X1 U2101 ( .IN1(AdderCntrl_ExcCheck_Datain[8]), .IN2(n1732), .OUT(n1989)
         );
  NAND3X1 U2102 ( .IN1(n1991), .IN2(n1990), .IN3(n1989), .OUT(n1992) );
  NOR2X1 U2103 ( .IN1(n1993), .IN2(n1992), .OUT(n2001) );
  NOR2X1 U2104 ( .IN1(MulCntrl_ExcCheck_Datain[9]), .IN2(
        MulCntrl_ExcCheck_Datain[8]), .OUT(n2000) );
  NOR2X1 U2105 ( .IN1(MulCntrl_ExcCheck_Datain[12]), .IN2(
        MulCntrl_ExcCheck_Datain[11]), .OUT(n1996) );
  NOR2X1 U2106 ( .IN1(MulCntrl_ExcCheck_Datain[14]), .IN2(
        MulCntrl_ExcCheck_Datain[13]), .OUT(n1995) );
  NOR2X1 U2107 ( .IN1(MulCntrl_ExcCheck_Datain[7]), .IN2(
        MulCntrl_ExcCheck_Datain[10]), .OUT(n1994) );
  NAND3X1 U2108 ( .IN1(n1996), .IN2(n1995), .IN3(n1994), .OUT(n1997) );
  NOR2X1 U2109 ( .IN1(n1998), .IN2(n1997), .OUT(n1999) );
  AOI22 U2110 ( .IN1(n2002), .IN2(n2001), .IN3(n2000), .IN4(n1999), .OUT(n2104) );
  OAI21 U2111 ( .IN1(n2106), .IN2(n2003), .IN3(n2104), .OUT(n2004) );
  OAI21 U2112 ( .IN1(n2107), .IN2(n1769), .IN3(n2005), .OUT(n1655) );
  OAI21 U2113 ( .IN1(n2107), .IN2(n1751), .IN3(n2005), .OUT(n1654) );
  AOI22 U2114 ( .IN1(u_booth_Q1_reg), .IN2(n1736), .IN3(n713), .IN4(n1743), 
        .OUT(n2021) );
  NOR2X1 U2115 ( .IN1(Booth_Add_ack), .IN2(n1868), .OUT(n2006) );
  NOR2X1 U2116 ( .IN1(u_Adder_interconnect_stateMC_1_), .IN2(n1739), .OUT(
        n2018) );
  NAND2X1 U2117 ( .IN1(Add_valid), .IN2(n1740), .OUT(n2007) );
  AOI22 U2118 ( .IN1(u_Adder_interconnect_stateMC_1_), .IN2(n1749), .IN3(n2018), .IN4(n2007), .OUT(n2009) );
  NAND3X1 U2119 ( .IN1(n1794), .IN2(u_Adder_interconnect_stateMC_1_), .IN3(
        n1739), .OUT(n2011) );
  OAI21 U2120 ( .IN1(n2009), .IN2(n2008), .IN3(n2011), .OUT(n1622) );
  NAND2X1 U2121 ( .IN1(Booth_Add_valid), .IN2(
        u_Adder_interconnect_priority_reg), .OUT(n2010) );
  AOI22 U2122 ( .IN1(n2018), .IN2(n2010), .IN3(n1739), .IN4(n1749), .OUT(n2013) );
  OAI21 U2123 ( .IN1(n2013), .IN2(n2012), .IN3(n2011), .OUT(n1621) );
  AOI22 U2124 ( .IN1(u_Adder_interconnect_priority_reg), .IN2(n1758), .IN3(
        Add_valid), .IN4(n1740), .OUT(n2015) );
  OAI21 U2125 ( .IN1(u_Adder_interconnect_priority_reg), .IN2(n2018), .IN3(
        n1794), .OUT(n2014) );
  AOI21 U2126 ( .IN1(n2018), .IN2(n2015), .IN3(n2014), .OUT(n1620) );
  NOR2X1 U2127 ( .IN1(n802), .IN2(u_adder_24b_StateMC_1_), .OUT(n2037) );
  NOR2X1 U2128 ( .IN1(n2037), .IN2(n2016), .OUT(n1589) );
  AOI21 U2129 ( .IN1(u_adder_24b_StateMC_1_), .IN2(n1770), .IN3(n2037), .OUT(
        n2017) );
  NOR2X1 U2130 ( .IN1(n2017), .IN2(n1795), .OUT(n1588) );
  NOR2X1 U2131 ( .IN1(n2018), .IN2(n1795), .OUT(n2095) );
  NOR2X1 U2132 ( .IN1(n1795), .IN2(n1749), .OUT(n2096) );
  AOI22 U2133 ( .IN1(Booth_Add_ack), .IN2(n2095), .IN3(n2019), .IN4(n2096), 
        .OUT(n2020) );
  AOI22 U2134 ( .IN1(n1867), .IN2(n1774), .IN3(n1866), .IN4(Add_dataout[6]), 
        .OUT(n2023) );
  AOI22 U2135 ( .IN1(n1867), .IN2(u_booth_A_reg_7_), .IN3(n1866), .IN4(
        Add_dataout[7]), .OUT(n2025) );
  AOI21 U2136 ( .IN1(n1746), .IN2(n584), .IN3(n1738), .OUT(n2027) );
  NAND2X1 U2137 ( .IN1(n1794), .IN2(n2027), .OUT(n2028) );
  OAI21 U2138 ( .IN1(n2029), .IN2(n2181), .IN3(n2028), .OUT(n1513) );
  AOI21 U2139 ( .IN1(n2182), .IN2(n2030), .IN3(MulCntrl_valid), .OUT(n2031) );
  OAI21 U2140 ( .IN1(n1738), .IN2(n1746), .IN3(n2031), .OUT(n2032) );
  NAND2X1 U2141 ( .IN1(n1794), .IN2(n2032), .OUT(n992) );
  AOI21 U2142 ( .IN1(n2034), .IN2(n2094), .IN3(n2033), .OUT(
        u_Adder_interconnect_N53) );
  AOI21 U2143 ( .IN1(n2036), .IN2(n2099), .IN3(n2035), .OUT(
        u_ExcChecker_interconnect_N53) );
  NAND3X1 U2144 ( .IN1(n1794), .IN2(n2037), .IN3(n768), .OUT(n2038) );
  NOR2X1 U2145 ( .IN1(n1771), .IN2(n2069), .OUT(n707) );
  NAND2X1 U2146 ( .IN1(n1737), .IN2(n1742), .OUT(n2062) );
  NOR2X1 U2147 ( .IN1(u_booth_M_reg_2_), .IN2(n2062), .OUT(n2057) );
  NOR2X1 U2148 ( .IN1(n2058), .IN2(u_booth_M_reg_3_), .OUT(n2053) );
  NOR2X1 U2149 ( .IN1(u_booth_M_reg_4_), .IN2(n2054), .OUT(n2049) );
  NOR2X1 U2150 ( .IN1(n2050), .IN2(u_booth_M_reg_5_), .OUT(n2045) );
  NOR2X1 U2151 ( .IN1(u_booth_M_reg_6_), .IN2(n2046), .OUT(n2041) );
  NOR2X1 U2152 ( .IN1(u_booth_Q1_reg), .IN2(n713), .OUT(n2039) );
  AOI21 U2153 ( .IN1(n2041), .IN2(n1750), .IN3(n2044), .OUT(n705) );
  NAND3X1 U2154 ( .IN1(u_booth_Q1_reg), .IN2(n713), .IN3(n2040), .OUT(n2043)
         );
  OAI21 U2155 ( .IN1(n1750), .IN2(n2041), .IN3(n705), .OUT(n2042) );
  OAI21 U2156 ( .IN1(n2043), .IN2(n1750), .IN3(n2042), .OUT(n704) );
  MUX2X1 U2157 ( .IN1(n2046), .IN2(n2045), .S(u_booth_M_reg_6_), .OUT(n2047)
         );
  AOI22 U2158 ( .IN1(u_booth_M_reg_6_), .IN2(n2065), .IN3(n2066), .IN4(n2047), 
        .OUT(n2048) );
  MUX2X1 U2159 ( .IN1(n2050), .IN2(n2049), .S(u_booth_M_reg_5_), .OUT(n2051)
         );
  AOI22 U2160 ( .IN1(u_booth_M_reg_5_), .IN2(n2065), .IN3(n2066), .IN4(n2051), 
        .OUT(n2052) );
  MUX2X1 U2161 ( .IN1(n2054), .IN2(n2053), .S(u_booth_M_reg_4_), .OUT(n2055)
         );
  AOI22 U2162 ( .IN1(u_booth_M_reg_4_), .IN2(n2065), .IN3(n2066), .IN4(n2055), 
        .OUT(n2056) );
  MUX2X1 U2163 ( .IN1(n2058), .IN2(n2057), .S(u_booth_M_reg_3_), .OUT(n2059)
         );
  AOI22 U2164 ( .IN1(u_booth_M_reg_3_), .IN2(n2065), .IN3(n2066), .IN4(n2059), 
        .OUT(n2060) );
  MUX2X1 U2165 ( .IN1(n2062), .IN2(n2061), .S(u_booth_M_reg_2_), .OUT(n2063)
         );
  AOI22 U2166 ( .IN1(u_booth_M_reg_2_), .IN2(n2065), .IN3(n2066), .IN4(n2063), 
        .OUT(n2064) );
  AOI21 U2167 ( .IN1(n2066), .IN2(n1737), .IN3(n2065), .OUT(n2068) );
  NAND2X1 U2168 ( .IN1(n2066), .IN2(u_booth_N258), .OUT(n2067) );
  AOI22 U2169 ( .IN1(u_booth_M_reg_1_), .IN2(n2068), .IN3(n2067), .IN4(n1742), 
        .OUT(n698) );
  NOR2X1 U2170 ( .IN1(n1737), .IN2(n2069), .OUT(n697) );
  OAI21 U2171 ( .IN1(n654), .IN2(n2071), .IN3(n2070), .OUT(n622) );
  AOI22 U2172 ( .IN1(u_booth_M_reg_7_), .IN2(n2081), .IN3(n2080), .IN4(
        Booth_datain1[7]), .OUT(n2073) );
  AOI22 U2173 ( .IN1(u_booth_M_reg_6_), .IN2(n2081), .IN3(n2080), .IN4(
        Booth_datain1[6]), .OUT(n2074) );
  AOI22 U2174 ( .IN1(u_booth_M_reg_5_), .IN2(n2081), .IN3(n2080), .IN4(
        Booth_datain1[5]), .OUT(n2075) );
  AOI22 U2175 ( .IN1(u_booth_M_reg_4_), .IN2(n2081), .IN3(n2080), .IN4(
        Booth_datain1[4]), .OUT(n2076) );
  AOI22 U2176 ( .IN1(u_booth_M_reg_3_), .IN2(n2081), .IN3(n2080), .IN4(
        Booth_datain1[3]), .OUT(n2077) );
  AOI22 U2177 ( .IN1(u_booth_M_reg_2_), .IN2(n2081), .IN3(n2080), .IN4(
        Booth_datain1[2]), .OUT(n2078) );
  AOI22 U2178 ( .IN1(u_booth_M_reg_1_), .IN2(n2081), .IN3(n2080), .IN4(
        Booth_datain1[1]), .OUT(n2079) );
  AOI22 U2179 ( .IN1(u_booth_N258), .IN2(n2081), .IN3(n2080), .IN4(
        Booth_datain1[0]), .OUT(n2082) );
  AOI21 U2180 ( .IN1(n768), .IN2(n1757), .IN3(n1795), .OUT(n2092) );
  AOI22 U2181 ( .IN1(Add_dataout[1]), .IN2(n1787), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N123), .OUT(n2083) );
  AOI22 U2182 ( .IN1(Add_dataout[2]), .IN2(n1787), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N124), .OUT(n2084) );
  AOI22 U2183 ( .IN1(Add_dataout[3]), .IN2(n1787), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N125), .OUT(n2085) );
  AOI22 U2184 ( .IN1(Add_dataout[4]), .IN2(n1787), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N126), .OUT(n2086) );
  AOI22 U2185 ( .IN1(Add_dataout[5]), .IN2(n1787), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N127), .OUT(n2087) );
  AOI22 U2186 ( .IN1(Add_dataout[6]), .IN2(n1787), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N128), .OUT(n2088) );
  AOI22 U2187 ( .IN1(Add_dataout[7]), .IN2(n1787), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N129), .OUT(n2089) );
  INVX1 U2188 ( .IN(n2089), .OUT(n599) );
  AOI22 U2189 ( .IN1(Add_dataout[8]), .IN2(n1787), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N130), .OUT(n2090) );
  INVX1 U2190 ( .IN(n2090), .OUT(n598) );
  AOI22 U2191 ( .IN1(u_adder_24b_N52), .IN2(u_adder_24b_N131), .IN3(n1787), 
        .IN4(Add_carryout), .OUT(n2091) );
  AOI22 U2192 ( .IN1(Add_dataout[0]), .IN2(n1787), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N122), .OUT(n2093) );
  AOI22 U2193 ( .IN1(n2097), .IN2(n2096), .IN3(n2095), .IN4(Add_ack), .OUT(
        n2098) );
  AOI22 U2194 ( .IN1(n2102), .IN2(AdderCntrl_Exc_Ack), .IN3(n2101), .IN4(n2100), .OUT(n2103) );
  OAI21 U2195 ( .IN1(n2106), .IN2(n2105), .IN3(n2104), .OUT(n2109) );
  AOI22 U2196 ( .IN1(u_exc_check_N45), .IN2(n2109), .IN3(n2108), .IN4(
        ExcCheck_value[2]), .OUT(n2110) );
  NOR2X1 U2197 ( .IN1(n2111), .IN2(n1795), .OUT(n2144) );
  NOR2X1 U2198 ( .IN1(n1791), .IN2(n1795), .OUT(n2143) );
  AOI22 U2199 ( .IN1(DIN2[0]), .IN2(n1790), .IN3(n1791), .IN4(MulCntrl_Op2[0]), 
        .OUT(n2112) );
  AOI22 U2200 ( .IN1(n1791), .IN2(MulCntrl_Op2[1]), .IN3(n1790), .IN4(DIN2[1]), 
        .OUT(n2113) );
  AOI22 U2201 ( .IN1(n1791), .IN2(MulCntrl_Op2[2]), .IN3(n1790), .IN4(DIN2[2]), 
        .OUT(n2114) );
  AOI22 U2202 ( .IN1(n1791), .IN2(MulCntrl_Op2[3]), .IN3(n1790), .IN4(DIN2[3]), 
        .OUT(n2115) );
  AOI22 U2203 ( .IN1(n2144), .IN2(MulCntrl_Op2[4]), .IN3(n1790), .IN4(DIN2[4]), 
        .OUT(n2116) );
  AOI22 U2204 ( .IN1(n2144), .IN2(MulCntrl_Op2[5]), .IN3(n1790), .IN4(DIN2[5]), 
        .OUT(n2117) );
  AOI22 U2205 ( .IN1(n2144), .IN2(MulCntrl_Op2[6]), .IN3(n1790), .IN4(DIN2[6]), 
        .OUT(n2118) );
  AOI22 U2206 ( .IN1(n1791), .IN2(MulCntrl_Op2[7]), .IN3(n1790), .IN4(DIN2[7]), 
        .OUT(n2119) );
  AOI22 U2207 ( .IN1(n1791), .IN2(MulCntrl_Op2[8]), .IN3(n1790), .IN4(DIN2[8]), 
        .OUT(n2120) );
  AOI22 U2208 ( .IN1(n1791), .IN2(MulCntrl_Op2[9]), .IN3(n1790), .IN4(DIN2[9]), 
        .OUT(n2121) );
  AOI22 U2209 ( .IN1(n1791), .IN2(MulCntrl_Op2[10]), .IN3(n1790), .IN4(
        DIN2[10]), .OUT(n2122) );
  AOI22 U2210 ( .IN1(n1791), .IN2(MulCntrl_Op2[11]), .IN3(n1790), .IN4(
        DIN2[11]), .OUT(n2123) );
  AOI22 U2211 ( .IN1(n1791), .IN2(MulCntrl_Op2[12]), .IN3(n1790), .IN4(
        DIN2[12]), .OUT(n2124) );
  AOI22 U2212 ( .IN1(n1791), .IN2(MulCntrl_Op2[13]), .IN3(n1790), .IN4(
        DIN2[13]), .OUT(n2125) );
  AOI22 U2213 ( .IN1(n1791), .IN2(MulCntrl_Op2[14]), .IN3(n1790), .IN4(
        DIN2[14]), .OUT(n2126) );
  AOI22 U2214 ( .IN1(n2144), .IN2(MulCntrl_Op2[15]), .IN3(n2143), .IN4(
        DIN2[15]), .OUT(n2127) );
  AOI22 U2215 ( .IN1(n2144), .IN2(MulCntrl_Op1[0]), .IN3(n2143), .IN4(DIN1[0]), 
        .OUT(n2128) );
  AOI22 U2216 ( .IN1(n2144), .IN2(MulCntrl_Op1[1]), .IN3(n2143), .IN4(DIN1[1]), 
        .OUT(n2129) );
  AOI22 U2217 ( .IN1(n2144), .IN2(MulCntrl_Op1[2]), .IN3(n2143), .IN4(DIN1[2]), 
        .OUT(n2130) );
  AOI22 U2218 ( .IN1(n1791), .IN2(MulCntrl_Op1[3]), .IN3(n1790), .IN4(DIN1[3]), 
        .OUT(n2131) );
  AOI22 U2219 ( .IN1(n1791), .IN2(MulCntrl_Op1[4]), .IN3(n1790), .IN4(DIN1[4]), 
        .OUT(n2132) );
  AOI22 U2220 ( .IN1(n1791), .IN2(MulCntrl_Op1[5]), .IN3(n1790), .IN4(DIN1[5]), 
        .OUT(n2133) );
  AOI22 U2221 ( .IN1(n1791), .IN2(MulCntrl_Op1[6]), .IN3(n1790), .IN4(DIN1[6]), 
        .OUT(n2134) );
  AOI22 U2222 ( .IN1(n1791), .IN2(n1733), .IN3(n1790), .IN4(DIN1[7]), .OUT(
        n2135) );
  AOI22 U2223 ( .IN1(n1791), .IN2(MulCntrl_Op1[8]), .IN3(n2143), .IN4(DIN1[8]), 
        .OUT(n2136) );
  AOI22 U2224 ( .IN1(n1791), .IN2(MulCntrl_Op1[9]), .IN3(n1790), .IN4(DIN1[9]), 
        .OUT(n2137) );
  AOI22 U2225 ( .IN1(n1791), .IN2(MulCntrl_Op1[10]), .IN3(n1790), .IN4(
        DIN1[10]), .OUT(n2138) );
  AOI22 U2226 ( .IN1(n1791), .IN2(MulCntrl_Op1[11]), .IN3(n2143), .IN4(
        DIN1[11]), .OUT(n2139) );
  AOI22 U2227 ( .IN1(n1791), .IN2(MulCntrl_Op1[12]), .IN3(n1790), .IN4(
        DIN1[12]), .OUT(n2140) );
  AOI22 U2228 ( .IN1(n1791), .IN2(MulCntrl_Op1[13]), .IN3(n1790), .IN4(
        DIN1[13]), .OUT(n2141) );
  AOI22 U2229 ( .IN1(n1791), .IN2(MulCntrl_Op1[14]), .IN3(n1790), .IN4(
        DIN1[14]), .OUT(n2142) );
  AOI22 U2230 ( .IN1(n2144), .IN2(MulCntrl_Op1[15]), .IN3(n1790), .IN4(
        DIN1[15]), .OUT(n2145) );
  NOR2X1 U2231 ( .IN1(n2146), .IN2(n1795), .OUT(n2178) );
  NOR2X1 U2232 ( .IN1(n1792), .IN2(n1795), .OUT(n2179) );
  AOI22 U2233 ( .IN1(DIN2[0]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op2[0]), .OUT(n2147) );
  AOI22 U2234 ( .IN1(DIN2[1]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op2[1]), .OUT(n2148) );
  AOI22 U2235 ( .IN1(DIN2[2]), .IN2(n2179), .IN3(n1792), .IN4(
        AdderCntrl_Op2[2]), .OUT(n2149) );
  AOI22 U2236 ( .IN1(DIN2[3]), .IN2(n2179), .IN3(n1792), .IN4(
        AdderCntrl_Op2[3]), .OUT(n2150) );
  AOI22 U2237 ( .IN1(DIN2[4]), .IN2(n2179), .IN3(n1792), .IN4(
        AdderCntrl_Op2[4]), .OUT(n2151) );
  AOI22 U2238 ( .IN1(DIN2[5]), .IN2(n2179), .IN3(n1792), .IN4(
        AdderCntrl_Op2[5]), .OUT(n2152) );
  AOI22 U2239 ( .IN1(DIN2[6]), .IN2(n2179), .IN3(n1792), .IN4(
        AdderCntrl_Op2[6]), .OUT(n2153) );
  AOI22 U2240 ( .IN1(DIN2[7]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op2[7]), .OUT(n2154) );
  AOI22 U2241 ( .IN1(DIN2[8]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op2[8]), .OUT(n2155) );
  AOI22 U2242 ( .IN1(DIN2[9]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op2[9]), .OUT(n2156) );
  AOI22 U2243 ( .IN1(DIN2[10]), .IN2(n2179), .IN3(n1792), .IN4(
        AdderCntrl_Op2[10]), .OUT(n2157) );
  AOI22 U2244 ( .IN1(DIN2[11]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op2[11]), .OUT(n2158) );
  AOI22 U2245 ( .IN1(DIN2[12]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op2[12]), .OUT(n2159) );
  AOI22 U2246 ( .IN1(DIN2[13]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op2[13]), .OUT(n2160) );
  AOI22 U2247 ( .IN1(DIN2[14]), .IN2(n1793), .IN3(n2178), .IN4(
        AdderCntrl_Op2[14]), .OUT(n2161) );
  AOI22 U2248 ( .IN1(DIN2[15]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op2[15]), .OUT(n2162) );
  AOI22 U2249 ( .IN1(DIN1[0]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op1[0]), .OUT(n2163) );
  AOI22 U2250 ( .IN1(DIN1[1]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op1[1]), .OUT(n2164) );
  AOI22 U2251 ( .IN1(DIN1[2]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op1[2]), .OUT(n2165) );
  AOI22 U2252 ( .IN1(DIN1[3]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op1[3]), .OUT(n2166) );
  AOI22 U2253 ( .IN1(DIN1[4]), .IN2(n1793), .IN3(n2178), .IN4(
        AdderCntrl_Op1[4]), .OUT(n2167) );
  AOI22 U2254 ( .IN1(DIN1[5]), .IN2(n1793), .IN3(n2178), .IN4(
        AdderCntrl_Op1[5]), .OUT(n2168) );
  AOI22 U2255 ( .IN1(DIN1[6]), .IN2(n1793), .IN3(n2178), .IN4(
        AdderCntrl_Op1[6]), .OUT(n2169) );
  AOI22 U2256 ( .IN1(DIN1[7]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op1[7]), .OUT(n2170) );
  AOI22 U2257 ( .IN1(DIN1[8]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op1[8]), .OUT(n2171) );
  AOI22 U2258 ( .IN1(DIN1[9]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op1[9]), .OUT(n2172) );
  AOI22 U2259 ( .IN1(DIN1[10]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op1[10]), .OUT(n2173) );
  AOI22 U2260 ( .IN1(DIN1[11]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op1[11]), .OUT(n2174) );
  AOI22 U2261 ( .IN1(DIN1[12]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op1[12]), .OUT(n2175) );
  AOI22 U2262 ( .IN1(DIN1[13]), .IN2(n1793), .IN3(n1792), .IN4(
        AdderCntrl_Op1[13]), .OUT(n2176) );
  AOI22 U2263 ( .IN1(DIN1[14]), .IN2(n1793), .IN3(n2178), .IN4(
        AdderCntrl_Op1[14]), .OUT(n2177) );
  AOI22 U2264 ( .IN1(DIN1[15]), .IN2(n1793), .IN3(n2178), .IN4(
        AdderCntrl_Op1[15]), .OUT(n2180) );
  AOI21 U2265 ( .IN1(n2182), .IN2(MulCntrl_Dataout_valid), .IN3(n1795), .OUT(
        n2201) );
  AOI22 U2266 ( .IN1(n2202), .IN2(MulCntrl_Dataout[15]), .IN3(n1788), .IN4(
        MultResult_reg[15]), .OUT(n2183) );
  AOI22 U2267 ( .IN1(n2202), .IN2(MulCntrl_Dataout[14]), .IN3(n1788), .IN4(
        MultResult_reg[14]), .OUT(n2184) );
  AOI22 U2268 ( .IN1(n2202), .IN2(MulCntrl_Dataout[13]), .IN3(n1788), .IN4(
        MultResult_reg[13]), .OUT(n2185) );
  AOI22 U2269 ( .IN1(n2202), .IN2(MulCntrl_Dataout[12]), .IN3(n1788), .IN4(
        MultResult_reg[12]), .OUT(n2186) );
  AOI22 U2270 ( .IN1(n2202), .IN2(MulCntrl_Dataout[11]), .IN3(n1788), .IN4(
        MultResult_reg[11]), .OUT(n2187) );
  AOI22 U2271 ( .IN1(n2202), .IN2(MulCntrl_Dataout[10]), .IN3(n1788), .IN4(
        MultResult_reg[10]), .OUT(n2188) );
  AOI22 U2272 ( .IN1(n2202), .IN2(MulCntrl_Dataout[9]), .IN3(n1788), .IN4(
        MultResult_reg[9]), .OUT(n2189) );
  AOI22 U2273 ( .IN1(n2202), .IN2(MulCntrl_Dataout[8]), .IN3(n1788), .IN4(
        MultResult_reg[8]), .OUT(n2190) );
  AOI22 U2274 ( .IN1(n2202), .IN2(MulCntrl_Dataout[7]), .IN3(n1788), .IN4(
        MultResult_reg[7]), .OUT(n2191) );
  AOI22 U2275 ( .IN1(n2202), .IN2(MulCntrl_Dataout[6]), .IN3(n1788), .IN4(
        MultResult_reg[6]), .OUT(n2192) );
  AOI22 U2276 ( .IN1(n2202), .IN2(MulCntrl_Dataout[5]), .IN3(n1788), .IN4(
        MultResult_reg[5]), .OUT(n2193) );
  AOI22 U2277 ( .IN1(n2202), .IN2(MulCntrl_Dataout[4]), .IN3(n1788), .IN4(
        MultResult_reg[4]), .OUT(n2194) );
  AOI22 U2278 ( .IN1(n2202), .IN2(MulCntrl_Dataout[3]), .IN3(n1788), .IN4(
        MultResult_reg[3]), .OUT(n2195) );
  AOI22 U2279 ( .IN1(n2202), .IN2(MulCntrl_Dataout[2]), .IN3(n1788), .IN4(
        MultResult_reg[2]), .OUT(n2196) );
  AOI22 U2280 ( .IN1(n2202), .IN2(MulCntrl_Dataout[1]), .IN3(n1788), .IN4(
        MultResult_reg[1]), .OUT(n2197) );
  AOI22 U2281 ( .IN1(n2202), .IN2(MulCntrl_Dataout[0]), .IN3(n1788), .IN4(
        MultResult_reg[0]), .OUT(n2198) );
  AOI22 U2282 ( .IN1(n2202), .IN2(MulCntrl_Exc[2]), .IN3(n1788), .IN4(
        MultExc_reg[2]), .OUT(n2199) );
  AOI22 U2283 ( .IN1(n2202), .IN2(MulCntrl_Exc[1]), .IN3(n1788), .IN4(
        MultExc_reg[1]), .OUT(n2200) );
  AOI22 U2284 ( .IN1(n2202), .IN2(MulCntrl_Exc[0]), .IN3(n1788), .IN4(
        MultExc_reg[0]), .OUT(n2203) );
  NOR2X1 U2285 ( .IN1(n2205), .IN2(n1795), .OUT(n2224) );
  AOI22 U2286 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[15]), .IN3(n1789), .IN4(
        AdderResult_reg[15]), .OUT(n2206) );
  AOI22 U2287 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[14]), .IN3(n1789), .IN4(
        AdderResult_reg[14]), .OUT(n2207) );
  AOI22 U2288 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[13]), .IN3(n1789), .IN4(
        AdderResult_reg[13]), .OUT(n2208) );
  AOI22 U2289 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[12]), .IN3(n1789), .IN4(
        AdderResult_reg[12]), .OUT(n2209) );
  AOI22 U2290 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[11]), .IN3(n1789), .IN4(
        AdderResult_reg[11]), .OUT(n2210) );
  AOI22 U2291 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[10]), .IN3(n1789), .IN4(
        AdderResult_reg[10]), .OUT(n2211) );
  AOI22 U2292 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[9]), .IN3(n1789), .IN4(
        AdderResult_reg[9]), .OUT(n2212) );
  AOI22 U2293 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[8]), .IN3(n1789), .IN4(
        AdderResult_reg[8]), .OUT(n2213) );
  AOI22 U2294 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[7]), .IN3(n1789), .IN4(
        AdderResult_reg[7]), .OUT(n2214) );
  AOI22 U2295 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[6]), .IN3(n1789), .IN4(
        AdderResult_reg[6]), .OUT(n2215) );
  AOI22 U2296 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[5]), .IN3(n1789), .IN4(
        AdderResult_reg[5]), .OUT(n2216) );
  AOI22 U2297 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[4]), .IN3(n1789), .IN4(
        AdderResult_reg[4]), .OUT(n2217) );
  AOI22 U2298 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[3]), .IN3(n1789), .IN4(
        AdderResult_reg[3]), .OUT(n2218) );
  AOI22 U2299 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[2]), .IN3(n1789), .IN4(
        AdderResult_reg[2]), .OUT(n2219) );
  AOI22 U2300 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[1]), .IN3(n1789), .IN4(
        AdderResult_reg[1]), .OUT(n2220) );
  AOI22 U2301 ( .IN1(n2225), .IN2(AdderCntrl_Dataout[0]), .IN3(n1789), .IN4(
        AdderResult_reg[0]), .OUT(n2221) );
  AOI22 U2302 ( .IN1(n2225), .IN2(AdderCntrl_Exc[2]), .IN3(n1789), .IN4(
        AddExc_reg[2]), .OUT(n2222) );
  AOI22 U2303 ( .IN1(n2225), .IN2(AdderCntrl_Exc[1]), .IN3(n1789), .IN4(
        AddExc_reg[1]), .OUT(n2223) );
  AOI22 U2304 ( .IN1(n2225), .IN2(AdderCntrl_Exc[0]), .IN3(n1789), .IN4(
        AddExc_reg[0]), .OUT(n2226) );
endmodule

