
module Adder_cntrl ( CLK, Datain1, Datain2, Data_valid, Dataout, Dataout_valid, 
        Exc, Mode, Debug, Adder_datain1, Adder_datain2, Adder_valid, 
        Adder_dataout, Adder_carryout, Adder_ack, ExcCheck_valid, Exc_value, 
        Exc_Ack, RSTn_BAR, ExcCheck_Datain_15_, ExcCheck_Datain_14_, 
        ExcCheck_Datain_13__BAR, ExcCheck_Datain_12_, ExcCheck_Datain_11_, 
        ExcCheck_Datain_9_, ExcCheck_Datain_8_, ExcCheck_Datain_6_, 
        ExcCheck_Datain_5_, ExcCheck_Datain_4_, ExcCheck_Datain_3_, 
        ExcCheck_Datain_2_, ExcCheck_Datain_1_, ExcCheck_Datain_0_, 
        ExcCheck_Datain_10__BAR, ExcCheck_Datain_7__BAR );
  input [15:0] Datain1;
  input [15:0] Datain2;
  output [15:0] Dataout;
  output [2:0] Exc;
  input [2:0] Mode;
  output [4:0] Debug;
  output [8:0] Adder_datain1;
  output [8:0] Adder_datain2;
  input [8:0] Adder_dataout;
  input [2:0] Exc_value;
  input CLK, Data_valid, Adder_carryout, Adder_ack, Exc_Ack, RSTn_BAR;
  output Dataout_valid, Adder_valid, ExcCheck_valid, ExcCheck_Datain_15_,
         ExcCheck_Datain_14_, ExcCheck_Datain_13__BAR, ExcCheck_Datain_12_,
         ExcCheck_Datain_11_, ExcCheck_Datain_9_, ExcCheck_Datain_8_,
         ExcCheck_Datain_6_, ExcCheck_Datain_5_, ExcCheck_Datain_4_,
         ExcCheck_Datain_3_, ExcCheck_Datain_2_, ExcCheck_Datain_1_,
         ExcCheck_Datain_0_, ExcCheck_Datain_10__BAR, ExcCheck_Datain_7__BAR;
  wire   N143, N144, N145, N146, N147, N148, N149, N150, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N164, N165, N166,
         Debug_valid_reg, Op1_Sign_reg, Op2_Sign_reg, Op2_Mantissa_reg_7_,
         exc_reg_0_, carry_reg, N252, N253, N254, N255, N256, N257, N258, N259,
         N270, N363, N364, N365, N366, N367, N368, N369, N376, N384, N392,
         N419, N420, N421, N422, N423, N424, N425, N430, N437, N445, N691,
         C405_DATA2_3, C405_DATA2_5, C405_DATA2_6, C405_DATA2_7, n73, n103,
         n109, n110, n111, n112, n113, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n212, n213, n214, n215, n216, n217, n218, n219,
         n222, n223, n274, n277, n664, n672, n915, n922, n991, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, add_x_35_A_9_, add_x_35_A_8_, add_x_35_A_7_,
         add_x_35_A_6_, add_x_35_A_5_, add_x_35_A_4_, add_x_35_A_3_,
         add_x_35_A_2_, add_x_35_A_1_, add_x_35_A_0_, C1_Z_3, C1_Z_2, C1_Z_1,
         C1_Z_0, C2_Z_0, DP_OP_982J1_125_6202_n102, DP_OP_982J1_125_6202_n101,
         DP_OP_982J1_125_6202_n100, DP_OP_982J1_125_6202_n97,
         DP_OP_982J1_125_6202_n91, DP_OP_982J1_125_6202_n72,
         DP_OP_982J1_125_6202_n55, DP_OP_982J1_125_6202_n54,
         DP_OP_982J1_125_6202_n53, DP_OP_982J1_125_6202_n52,
         DP_OP_982J1_125_6202_n51, DP_OP_982J1_125_6202_n50,
         DP_OP_982J1_125_6202_n49, DP_OP_981J1_124_6202_n55,
         DP_OP_981J1_124_6202_n54, DP_OP_981J1_124_6202_n53,
         DP_OP_981J1_124_6202_n52, DP_OP_981J1_124_6202_n51,
         DP_OP_981J1_124_6202_n50, DP_OP_981J1_124_6202_n49,
         DP_OP_986_157_3518_n93, DP_OP_986_157_3518_n76,
         DP_OP_986_157_3518_n72, DP_OP_986_157_3518_n70,
         DP_OP_986_157_3518_n68, DP_OP_986_157_3518_n66,
         DP_OP_986_157_3518_n65, DP_OP_986_157_3518_n64,
         DP_OP_986_157_3518_n62, DP_OP_986_157_3518_n61,
         DP_OP_986_157_3518_n56, DP_OP_986_157_3518_n54,
         DP_OP_986_157_3518_n53, DP_OP_986_157_3518_n52,
         DP_OP_986_157_3518_n51, DP_OP_986_157_3518_n50,
         DP_OP_986_157_3518_n49, DP_OP_986_157_3518_n45,
         DP_OP_986_157_3518_n43, DP_OP_986_157_3518_n42,
         DP_OP_986_157_3518_n41, DP_OP_986_157_3518_n40,
         DP_OP_986_157_3518_n38, DP_OP_986_157_3518_n37,
         DP_OP_986_157_3518_n36, DP_OP_986_157_3518_n35,
         DP_OP_986_157_3518_n34, DP_OP_986_157_3518_n33,
         DP_OP_986_157_3518_n32, DP_OP_986_157_3518_n30,
         DP_OP_986_157_3518_n29, DP_OP_986_157_3518_n28,
         DP_OP_986_157_3518_n24, DP_OP_986_157_3518_n12,
         DP_OP_986_157_3518_n11, DP_OP_986_157_3518_n7, DP_OP_986_157_3518_n2,
         DP_OP_986_157_3518_n1, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n104, n105, n106, n107, n108, n114,
         n115, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n220, n221, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n275, n276, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n665, n666, n667, n668, n669, n670, n671, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n781, n782, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n916, n917, n918, n919, n920, n921,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203;
  wire   [2:0] StateMC;
  wire   [3:0] Debug_reg;
  wire   [7:0] Final_Exponent_reg;
  wire   [10:1] Final_Mantissa_reg;

  DFFRX1 Add_sign_reg_reg ( .D(n1103), .CLK(CLK), .CLRB(n73), .Q(n230), .QB(
        n277) );
  DFFRX1 Final_Mantissa_reg_reg_10_ ( .D(n1062), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[10]), .QB(n205) );
  DFFRX1 Final_Exponent_reg_reg_7_ ( .D(n1102), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[7]) );
  DFFRX1 StateMC_reg_1_ ( .D(n922), .CLK(CLK), .CLRB(n73), .Q(n220), .QB(
        StateMC[1]) );
  DFFRX1 Op2_Sign_reg_reg ( .D(n1090), .CLK(CLK), .CLRB(n73), .Q(Op2_Sign_reg), 
        .QB(n229) );
  DFFRX1 G_reg_reg ( .D(n1072), .CLK(CLK), .CLRB(n73), .Q(n226), .QB(
        add_x_35_A_2_) );
  DFFRX1 Final_Mantissa_reg_reg_2_ ( .D(n664), .CLK(CLK), .CLRB(n73), .Q(n208), 
        .QB(Final_Mantissa_reg[2]) );
  DFFRX1 Final_Mantissa_reg_reg_1_ ( .D(n672), .CLK(CLK), .CLRB(n73), .Q(n238), 
        .QB(Final_Mantissa_reg[1]) );
  DFFRX1 Final_Mantissa_reg_reg_0_ ( .D(n113), .CLK(CLK), .CLRB(n73), .Q(N691), 
        .QB(n236) );
  DFFRX1 Final_Mantissa_reg_reg_8_ ( .D(n1064), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[8]), .QB(n209) );
  DFFRX1 exc_reg_reg_0_ ( .D(n1092), .CLK(CLK), .CLRB(n73), .Q(exc_reg_0_), 
        .QB(n243) );
  DFFRX1 StateMC_reg_0_ ( .D(n991), .CLK(CLK), .CLRB(n73), .Q(n241), .QB(
        StateMC[0]) );
  DFFRX1 StateMC_reg_2_ ( .D(n915), .CLK(CLK), .CLRB(n73), .Q(n204), .QB(
        StateMC[2]) );
  DFFRX1 Op1_Sign_reg_reg ( .D(n1081), .CLK(CLK), .CLRB(n73), .Q(Op1_Sign_reg), 
        .QB(n228) );
  DFFRX1 Op1_Mantissa_reg_reg_6_ ( .D(n1083), .CLK(CLK), .CLRB(n73), .QB(n213)
         );
  DFFRX1 Op1_Mantissa_reg_reg_5_ ( .D(n1084), .CLK(CLK), .CLRB(n73), .QB(n214)
         );
  DFFRX1 Op1_Mantissa_reg_reg_4_ ( .D(n1085), .CLK(CLK), .CLRB(n73), .QB(n215)
         );
  DFFRX1 Op1_Mantissa_reg_reg_3_ ( .D(n1086), .CLK(CLK), .CLRB(n73), .QB(n216)
         );
  DFFRX1 Op1_Mantissa_reg_reg_2_ ( .D(n1087), .CLK(CLK), .CLRB(n73), .QB(n217)
         );
  DFFRX1 Op1_Mantissa_reg_reg_1_ ( .D(n1088), .CLK(CLK), .CLRB(n73), .QB(n218)
         );
  DFFRX1 Op1_Mantissa_reg_reg_0_ ( .D(n1089), .CLK(CLK), .CLRB(n73), .QB(n219)
         );
  DFFRX1 Op2_Mantissa_reg_reg_7_ ( .D(n1073), .CLK(CLK), .CLRB(n73), .Q(
        Op2_Mantissa_reg_7_), .QB(n244) );
  DFFRX1 R_reg_reg ( .D(n1070), .CLK(CLK), .CLRB(n73), .Q(n240), .QB(
        add_x_35_A_1_) );
  DFFRX1 S_reg_reg ( .D(n1071), .CLK(CLK), .CLRB(n73), .Q(n211), .QB(
        add_x_35_A_0_) );
  DFFRX1 Adder_datain2_reg_8_ ( .D(n124), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[8]) );
  DFFRX1 Adder_datain2_reg_7_ ( .D(n123), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[7]) );
  DFFRX1 Adder_datain1_reg_6_ ( .D(N258), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[6]) );
  DFFRX1 Adder_datain1_reg_5_ ( .D(N257), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[5]) );
  DFFRX1 Adder_datain1_reg_4_ ( .D(N256), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[4]) );
  DFFRX1 Adder_datain1_reg_3_ ( .D(N255), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[3]) );
  DFFRX1 Adder_datain1_reg_2_ ( .D(N254), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[2]) );
  DFFRX1 Adder_datain1_reg_1_ ( .D(N253), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[1]) );
  DFFRX1 Adder_datain1_reg_0_ ( .D(N252), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[0]) );
  DFFRX1 carry_reg_reg ( .D(n1061), .CLK(CLK), .CLRB(n73), .Q(carry_reg), .QB(
        n227) );
  DFFRX1 Final_Mantissa_reg_reg_9_ ( .D(n1063), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[9]), .QB(n232) );
  DFFRX1 Final_Mantissa_reg_reg_7_ ( .D(n1065), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[7]), .QB(n231) );
  DFFRX1 Final_Mantissa_reg_reg_6_ ( .D(n1066), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[6]), .QB(n206) );
  DFFRX1 Final_Mantissa_reg_reg_5_ ( .D(n1067), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[5]), .QB(n237) );
  DFFRX1 Final_Mantissa_reg_reg_4_ ( .D(n1068), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[4]), .QB(n233) );
  DFFRX1 Final_Mantissa_reg_reg_3_ ( .D(n1069), .CLK(CLK), .CLRB(n73), .Q(
        Final_Mantissa_reg[3]), .QB(n210) );
  DFFRX1 Debug_valid_reg_reg ( .D(n103), .CLK(CLK), .CLRB(n73), .Q(
        Debug_valid_reg), .QB(n246) );
  DFFRX1 Adder_valid_reg ( .D(n1091), .CLK(CLK), .CLRB(n73), .Q(Adder_valid), 
        .QB(n245) );
  DFFRX1 exc_reg_reg_1_ ( .D(n1093), .CLK(CLK), .CLRB(n73), .Q(n242), .QB(n223) );
  DFFRX1 exc_reg_reg_2_ ( .D(n1101), .CLK(CLK), .CLRB(n73), .QB(n222) );
  DFFRX1 Final_Sign_reg_reg ( .D(n1060), .CLK(CLK), .CLRB(n73), .Q(n251), .QB(
        n274) );
  DFFRX1 Op1_Mantissa_reg_reg_7_ ( .D(n1082), .CLK(CLK), .CLRB(n73), .QB(n212)
         );
  DFFRX1 Adder_datain1_reg_7_ ( .D(N259), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain1[7]) );
  DFFRX1 Op2_Mantissa_reg_reg_0_ ( .D(n1080), .CLK(CLK), .CLRB(n73), .Q(n250), 
        .QB(add_x_35_A_3_) );
  DFFRX1 Adder_datain2_reg_0_ ( .D(n116), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[0]) );
  DFFRX1 Op2_Mantissa_reg_reg_1_ ( .D(n1079), .CLK(CLK), .CLRB(n73), .Q(n225), 
        .QB(add_x_35_A_4_) );
  DFFRX1 Adder_datain2_reg_1_ ( .D(n117), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[1]) );
  DFFRX1 Op2_Mantissa_reg_reg_2_ ( .D(n1078), .CLK(CLK), .CLRB(n73), .Q(n249), 
        .QB(add_x_35_A_5_) );
  DFFRX1 Adder_datain2_reg_2_ ( .D(n118), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[2]) );
  DFFRX1 Op2_Mantissa_reg_reg_3_ ( .D(n1077), .CLK(CLK), .CLRB(n73), .Q(n221), 
        .QB(add_x_35_A_6_) );
  DFFRX1 Adder_datain2_reg_3_ ( .D(n119), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[3]) );
  DFFRX1 Op2_Mantissa_reg_reg_4_ ( .D(n1076), .CLK(CLK), .CLRB(n73), .Q(n248), 
        .QB(add_x_35_A_7_) );
  DFFRX1 Adder_datain2_reg_4_ ( .D(n120), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[4]) );
  DFFRX1 Op2_Mantissa_reg_reg_5_ ( .D(n1075), .CLK(CLK), .CLRB(n73), .Q(n224), 
        .QB(add_x_35_A_8_) );
  DFFRX1 Adder_datain2_reg_5_ ( .D(n121), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[5]) );
  DFFRX1 Op2_Mantissa_reg_reg_6_ ( .D(n1074), .CLK(CLK), .CLRB(n73), .Q(n247), 
        .QB(add_x_35_A_9_) );
  DFFRX1 Adder_datain2_reg_6_ ( .D(n122), .CLK(CLK), .CLRB(n73), .Q(
        Adder_datain2[6]) );
  DFFRX1 Final_Exponent_reg_reg_0_ ( .D(n1094), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[0]), .QB(n235) );
  DFFRX1 Final_Exponent_reg_reg_1_ ( .D(n1095), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[1]), .QB(n239) );
  DFFRX1 Final_Exponent_reg_reg_2_ ( .D(n1096), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[2]), .QB(n207) );
  DFFRX1 Final_Exponent_reg_reg_3_ ( .D(n1097), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[3]), .QB(n234) );
  DFFRX1 Final_Exponent_reg_reg_4_ ( .D(n1098), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[4]) );
  DFFRX1 Final_Exponent_reg_reg_5_ ( .D(n1099), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[5]) );
  DFFRX1 Final_Exponent_reg_reg_6_ ( .D(n1100), .CLK(CLK), .CLRB(n73), .Q(
        Final_Exponent_reg[6]), .QB(n155) );
  DFFRX1 ExcCheck_valid_reg ( .D(N270), .CLK(CLK), .CLRB(n73), .Q(
        ExcCheck_valid) );
  DFFRX1 Debug_reg_reg_3_ ( .D(n112), .CLK(CLK), .CLRB(n73), .Q(Debug_reg[3])
         );
  DFFRX1 Debug_reg_reg_2_ ( .D(n111), .CLK(CLK), .CLRB(n73), .Q(Debug_reg[2])
         );
  DFFRX1 Debug_reg_reg_1_ ( .D(n110), .CLK(CLK), .CLRB(n73), .Q(Debug_reg[1])
         );
  DFFRX1 Debug_reg_reg_0_ ( .D(n109), .CLK(CLK), .CLRB(n73), .Q(Debug_reg[0])
         );
  FULLADD DP_OP_982J1_125_6202_U62 ( .A(n194), .B(Datain2[8]), .CIN(
        DP_OP_982J1_125_6202_n55), .COUT(DP_OP_982J1_125_6202_n54), .SUM(N419)
         );
  FULLADD DP_OP_982J1_125_6202_U61 ( .A(n195), .B(DP_OP_982J1_125_6202_n97), 
        .CIN(DP_OP_982J1_125_6202_n54), .COUT(DP_OP_982J1_125_6202_n53), .SUM(
        N420) );
  FULLADD DP_OP_982J1_125_6202_U60 ( .A(n196), .B(Datain2[10]), .CIN(
        DP_OP_982J1_125_6202_n53), .COUT(DP_OP_982J1_125_6202_n52), .SUM(N421)
         );
  FULLADD DP_OP_982J1_125_6202_U59 ( .A(n198), .B(Datain2[11]), .CIN(
        DP_OP_982J1_125_6202_n52), .COUT(DP_OP_982J1_125_6202_n51), .SUM(N422)
         );
  FULLADD DP_OP_982J1_125_6202_U58 ( .A(n199), .B(DP_OP_982J1_125_6202_n100), 
        .CIN(DP_OP_982J1_125_6202_n51), .COUT(DP_OP_982J1_125_6202_n50), .SUM(
        N423) );
  FULLADD DP_OP_982J1_125_6202_U57 ( .A(n200), .B(DP_OP_982J1_125_6202_n101), 
        .CIN(DP_OP_982J1_125_6202_n50), .COUT(DP_OP_982J1_125_6202_n49), .SUM(
        N424) );
  FULLADD DP_OP_981J1_124_6202_U62 ( .A(n176), .B(Datain1[8]), .CIN(
        DP_OP_981J1_124_6202_n55), .COUT(DP_OP_981J1_124_6202_n54), .SUM(N363)
         );
  FULLADD DP_OP_981J1_124_6202_U61 ( .A(n177), .B(Datain1[9]), .CIN(
        DP_OP_981J1_124_6202_n54), .COUT(DP_OP_981J1_124_6202_n53), .SUM(N364)
         );
  FULLADD DP_OP_981J1_124_6202_U60 ( .A(n178), .B(Datain1[10]), .CIN(
        DP_OP_981J1_124_6202_n53), .COUT(DP_OP_981J1_124_6202_n52), .SUM(N365)
         );
  FULLADD DP_OP_981J1_124_6202_U59 ( .A(n179), .B(DP_OP_982J1_125_6202_n91), 
        .CIN(DP_OP_981J1_124_6202_n52), .COUT(DP_OP_981J1_124_6202_n51), .SUM(
        N366) );
  FULLADD DP_OP_981J1_124_6202_U58 ( .A(n144), .B(Datain1[12]), .CIN(
        DP_OP_981J1_124_6202_n51), .COUT(DP_OP_981J1_124_6202_n50), .SUM(N367)
         );
  NAND2X1 DP_OP_986_157_3518_U28 ( .IN1(DP_OP_986_157_3518_n53), .IN2(
        DP_OP_986_157_3518_n37), .OUT(DP_OP_986_157_3518_n24) );
  NAND2X1 DP_OP_986_157_3518_U23 ( .IN1(DP_OP_986_157_3518_n12), .IN2(
        DP_OP_986_157_3518_n11), .OUT(C405_DATA2_3) );
  NAND2X1 DP_OP_986_157_3518_U22 ( .IN1(C2_Z_0), .IN2(Final_Exponent_reg[4]), 
        .OUT(DP_OP_986_157_3518_n34) );
  NAND2X1 DP_OP_986_157_3518_U62 ( .IN1(C2_Z_0), .IN2(Final_Exponent_reg[0]), 
        .OUT(DP_OP_986_157_3518_n50) );
  NAND2X1 DP_OP_986_157_3518_U1 ( .IN1(DP_OP_986_157_3518_n2), .IN2(
        DP_OP_986_157_3518_n1), .OUT(C405_DATA2_7) );
  NANDX2 DP_OP_986_157_3518_U42 ( .IN1(DP_OP_986_157_3518_n68), .IN2(
        Final_Exponent_reg[2]), .OUT(DP_OP_986_157_3518_n42) );
  NANDX2 DP_OP_986_157_3518_U31 ( .IN1(DP_OP_986_157_3518_n64), .IN2(
        DP_OP_986_157_3518_n93), .OUT(DP_OP_986_157_3518_n37) );
  NANDX2 DP_OP_986_157_3518_U69 ( .IN1(DP_OP_986_157_3518_n66), .IN2(
        DP_OP_986_157_3518_n65), .OUT(DP_OP_986_157_3518_n68) );
  NANDX2 DP_OP_986_157_3518_U51 ( .IN1(DP_OP_986_157_3518_n72), .IN2(
        Final_Exponent_reg[1]), .OUT(DP_OP_986_157_3518_n45) );
  NANDX2 DP_OP_986_157_3518_U65 ( .IN1(DP_OP_986_157_3518_n62), .IN2(
        DP_OP_986_157_3518_n61), .OUT(DP_OP_986_157_3518_n64) );
  NOR2X1 DP_OP_986_157_3518_U61 ( .IN1(Final_Exponent_reg[0]), .IN2(C2_Z_0), 
        .OUT(DP_OP_986_157_3518_n49) );
  NOR2X1 DP_OP_986_157_3518_U41 ( .IN1(Final_Exponent_reg[2]), .IN2(
        DP_OP_986_157_3518_n68), .OUT(DP_OP_986_157_3518_n41) );
  AOI21 DP_OP_986_157_3518_U36 ( .IN1(DP_OP_986_157_3518_n43), .IN2(
        DP_OP_986_157_3518_n54), .IN3(DP_OP_986_157_3518_n40), .OUT(
        DP_OP_986_157_3518_n38) );
  NOR2X1 DP_OP_986_157_3518_U30 ( .IN1(DP_OP_986_157_3518_n93), .IN2(
        DP_OP_986_157_3518_n64), .OUT(DP_OP_986_157_3518_n36) );
  OAI21 DP_OP_986_157_3518_U27 ( .IN1(DP_OP_986_157_3518_n36), .IN2(
        DP_OP_986_157_3518_n38), .IN3(DP_OP_986_157_3518_n37), .OUT(
        DP_OP_986_157_3518_n35) );
  NOR2X1 DP_OP_986_157_3518_U21 ( .IN1(Final_Exponent_reg[4]), .IN2(C2_Z_0), 
        .OUT(DP_OP_986_157_3518_n33) );
  AOI21 DP_OP_986_157_3518_U16 ( .IN1(DP_OP_986_157_3518_n35), .IN2(
        DP_OP_986_157_3518_n52), .IN3(DP_OP_986_157_3518_n32), .OUT(
        DP_OP_986_157_3518_n30) );
  FULLADD DP_OP_986_157_3518_U10 ( .A(C2_Z_0), .B(n145), .CIN(
        DP_OP_986_157_3518_n51), .COUT(DP_OP_986_157_3518_n29), .SUM(
        C405_DATA2_5) );
  FULLADD DP_OP_986_157_3518_U9 ( .A(C2_Z_0), .B(n156), .CIN(
        DP_OP_986_157_3518_n29), .COUT(DP_OP_986_157_3518_n28), .SUM(
        C405_DATA2_6) );
  NOR2X1 U3 ( .IN1(n360), .IN2(n361), .OUT(n1) );
  NAND3X1 U4 ( .IN1(n602), .IN2(n362), .IN3(n1), .OUT(n373) );
  NAND3X1 U5 ( .IN1(n431), .IN2(n280), .IN3(n281), .OUT(n536) );
  AOI22 U6 ( .IN1(n156), .IN2(n647), .IN3(n822), .IN4(Datain1[13]), .OUT(n2)
         );
  NAND2X1 U7 ( .IN1(DP_OP_982J1_125_6202_n101), .IN2(n821), .OUT(n3) );
  NAND2X1 U8 ( .IN1(C405_DATA2_6), .IN2(n650), .OUT(n4) );
  NAND3X1 U9 ( .IN1(n2), .IN2(n3), .IN3(n4), .OUT(n1100) );
  INVX1 U10 ( .IN(n657), .OUT(n5) );
  AOI22 U11 ( .IN1(n691), .IN2(n772), .IN3(n666), .IN4(n5), .OUT(n6) );
  INVX1 U12 ( .IN(n663), .OUT(n7) );
  INVX1 U13 ( .IN(n662), .OUT(n8) );
  AOI22 U14 ( .IN1(n685), .IN2(n661), .IN3(n7), .IN4(n8), .OUT(n9) );
  AOI22 U15 ( .IN1(n659), .IN2(n671), .IN3(n752), .IN4(n674), .OUT(n10) );
  AOI22 U16 ( .IN1(n658), .IN2(n676), .IN3(n665), .IN4(n684), .OUT(n11) );
  NAND3X1 U17 ( .IN1(n9), .IN2(n10), .IN3(n11), .OUT(n12) );
  AOI21 U18 ( .IN1(n656), .IN2(n690), .IN3(n12), .OUT(n13) );
  NAND2X1 U19 ( .IN1(n6), .IN2(n13), .OUT(n706) );
  NAND3X1 U20 ( .IN1(n757), .IN2(n631), .IN3(n675), .OUT(n14) );
  INVX1 U21 ( .IN(n14), .OUT(n15) );
  NAND3X1 U22 ( .IN1(n594), .IN2(n694), .IN3(n15), .OUT(n718) );
  INVX1 U23 ( .IN(n820), .OUT(n16) );
  AOI21 U24 ( .IN1(n380), .IN2(n827), .IN3(n16), .OUT(n539) );
  AOI22 U25 ( .IN1(n145), .IN2(n647), .IN3(n822), .IN4(Datain1[12]), .OUT(n17)
         );
  NAND2X1 U26 ( .IN1(C405_DATA2_5), .IN2(n650), .OUT(n18) );
  NAND2X1 U27 ( .IN1(DP_OP_982J1_125_6202_n100), .IN2(n821), .OUT(n19) );
  NAND3X1 U28 ( .IN1(n17), .IN2(n19), .IN3(n18), .OUT(n1099) );
  INVX1 U29 ( .IN(n610), .OUT(n20) );
  OAI21 U30 ( .IN1(n609), .IN2(n20), .IN3(n643), .OUT(n617) );
  NAND3X1 U31 ( .IN1(n691), .IN2(n207), .IN3(n239), .OUT(n663) );
  NAND3X1 U32 ( .IN1(n204), .IN2(Adder_ack), .IN3(n726), .OUT(n1138) );
  NAND3X1 U33 ( .IN1(n608), .IN2(n316), .IN3(n618), .OUT(n21) );
  INVX1 U34 ( .IN(n21), .OUT(n22) );
  NAND3X1 U35 ( .IN1(n694), .IN2(n669), .IN3(n22), .OUT(n769) );
  INVX1 U36 ( .IN(n494), .OUT(n23) );
  NOR2X1 U37 ( .IN1(n466), .IN2(n23), .OUT(n554) );
  AOI22 U38 ( .IN1(Final_Exponent_reg[4]), .IN2(n647), .IN3(n822), .IN4(
        DP_OP_982J1_125_6202_n91), .OUT(n24) );
  INVX1 U39 ( .IN(DP_OP_986_157_3518_n35), .OUT(n25) );
  NAND2X1 U40 ( .IN1(DP_OP_986_157_3518_n34), .IN2(DP_OP_986_157_3518_n52), 
        .OUT(n26) );
  OAI21 U41 ( .IN1(n25), .IN2(n26), .IN3(n650), .OUT(n27) );
  AOI21 U42 ( .IN1(n25), .IN2(n26), .IN3(n27), .OUT(n28) );
  AOI21 U43 ( .IN1(n821), .IN2(Datain2[11]), .IN3(n28), .OUT(n29) );
  NAND2X1 U44 ( .IN1(n24), .IN2(n29), .OUT(n1098) );
  INVX1 U45 ( .IN(n815), .OUT(n30) );
  NOR2X1 U46 ( .IN1(n1134), .IN2(n30), .OUT(n31) );
  MUX2X1 U47 ( .IN1(add_x_35_A_6_), .IN2(n221), .S(n31), .OUT(n32) );
  NOR2X1 U48 ( .IN1(n1130), .IN2(n32), .OUT(n119) );
  OAI21 U49 ( .IN1(C1_Z_0), .IN2(C2_Z_0), .IN3(n163), .OUT(n33) );
  INVX4 U50 ( .IN(n33), .OUT(DP_OP_986_157_3518_n76) );
  INVX1 U51 ( .IN(n1000), .OUT(n34) );
  NAND3X1 U52 ( .IN1(n273), .IN2(n271), .IN3(n1120), .OUT(n35) );
  NAND2X1 U53 ( .IN1(N160), .IN2(n34), .OUT(n36) );
  AOI21 U54 ( .IN1(n35), .IN2(n36), .IN3(n1001), .OUT(n1016) );
  AOI22 U55 ( .IN1(Final_Exponent_reg[2]), .IN2(n647), .IN3(n822), .IN4(
        Datain1[9]), .OUT(n37) );
  NAND2X1 U56 ( .IN1(DP_OP_986_157_3518_n42), .IN2(DP_OP_986_157_3518_n54), 
        .OUT(n38) );
  INVX1 U57 ( .IN(DP_OP_986_157_3518_n43), .OUT(n39) );
  OAI21 U58 ( .IN1(n38), .IN2(n39), .IN3(n650), .OUT(n40) );
  AOI21 U59 ( .IN1(n38), .IN2(n39), .IN3(n40), .OUT(n41) );
  AOI21 U60 ( .IN1(n821), .IN2(DP_OP_982J1_125_6202_n97), .IN3(n41), .OUT(n42)
         );
  NAND2X1 U61 ( .IN1(n37), .IN2(n42), .OUT(n1096) );
  INVX1 U62 ( .IN(n815), .OUT(n43) );
  NOR2X1 U63 ( .IN1(n1136), .IN2(n43), .OUT(n44) );
  MUX2X1 U64 ( .IN1(add_x_35_A_4_), .IN2(n225), .S(n44), .OUT(n45) );
  NOR2X1 U65 ( .IN1(n1130), .IN2(n45), .OUT(n117) );
  OAI21 U66 ( .IN1(n279), .IN2(n395), .IN3(n402), .OUT(n46) );
  NOR2X1 U67 ( .IN1(n535), .IN2(n46), .OUT(n47) );
  AOI22 U68 ( .IN1(n279), .IN2(n546), .IN3(n276), .IN4(n473), .OUT(n48) );
  AOI22 U69 ( .IN1(n278), .IN2(n450), .IN3(n275), .IN4(n474), .OUT(n49) );
  AOI21 U70 ( .IN1(n48), .IN2(n49), .IN3(n516), .OUT(n50) );
  AOI22 U71 ( .IN1(n280), .IN2(n537), .IN3(n826), .IN4(Adder_dataout[3]), 
        .OUT(n51) );
  AOI22 U72 ( .IN1(n481), .IN2(n526), .IN3(n477), .IN4(n548), .OUT(n52) );
  NOR2X1 U73 ( .IN1(n47), .IN2(n50), .OUT(n53) );
  NAND3X1 U74 ( .IN1(n52), .IN2(n51), .IN3(n53), .OUT(n54) );
  AOI21 U75 ( .IN1(n439), .IN2(n528), .IN3(n54), .OUT(n55) );
  AOI22 U76 ( .IN1(n445), .IN2(n479), .IN3(n482), .IN4(n513), .OUT(n56) );
  AOI22 U77 ( .IN1(n481), .IN2(n484), .IN3(n486), .IN4(n456), .OUT(n57) );
  NAND2X1 U78 ( .IN1(n56), .IN2(n57), .OUT(n58) );
  AOI22 U79 ( .IN1(n279), .IN2(n518), .IN3(n487), .IN4(n58), .OUT(n59) );
  OAI21 U80 ( .IN1(RSTn_BAR), .IN2(n55), .IN3(n59), .OUT(n1066) );
  AOI22 U81 ( .IN1(n230), .IN2(carry_reg), .IN3(n227), .IN4(n277), .OUT(n60)
         );
  INVX1 U82 ( .IN(n60), .OUT(n328) );
  INVX1 U83 ( .IN(C2_Z_0), .OUT(n61) );
  INVX1 U84 ( .IN(Final_Exponent_reg[7]), .OUT(n62) );
  AOI22 U85 ( .IN1(Final_Exponent_reg[7]), .IN2(C2_Z_0), .IN3(n61), .IN4(n62), 
        .OUT(DP_OP_986_157_3518_n7) );
  INVX1 U86 ( .IN(Final_Mantissa_reg[10]), .OUT(n63) );
  OAI21 U87 ( .IN1(n338), .IN2(n63), .IN3(n353), .OUT(n360) );
  INVX1 U88 ( .IN(N159), .OUT(n64) );
  AOI22 U89 ( .IN1(N159), .IN2(Datain1[3]), .IN3(Datain1[2]), .IN4(n64), .OUT(
        n65) );
  AOI22 U90 ( .IN1(N159), .IN2(Datain1[1]), .IN3(Datain1[0]), .IN4(n64), .OUT(
        n66) );
  INVX1 U91 ( .IN(N160), .OUT(n67) );
  AOI22 U92 ( .IN1(N160), .IN2(n65), .IN3(n66), .IN4(n67), .OUT(n68) );
  AOI22 U93 ( .IN1(N159), .IN2(Datain1[7]), .IN3(Datain1[6]), .IN4(n64), .OUT(
        n69) );
  AOI22 U94 ( .IN1(N159), .IN2(n273), .IN3(Datain1[4]), .IN4(n64), .OUT(n70)
         );
  AOI22 U95 ( .IN1(N160), .IN2(n69), .IN3(n70), .IN4(n67), .OUT(n71) );
  MUX2X1 U96 ( .IN1(n68), .IN2(n71), .S(N161), .OUT(n1188) );
  AOI22 U97 ( .IN1(Final_Exponent_reg[1]), .IN2(n647), .IN3(n822), .IN4(
        Datain1[8]), .OUT(n72) );
  INVX1 U98 ( .IN(n165), .OUT(n74) );
  NAND2X1 U99 ( .IN1(DP_OP_986_157_3518_n45), .IN2(n168), .OUT(n75) );
  OAI21 U100 ( .IN1(n74), .IN2(n75), .IN3(n650), .OUT(n76) );
  AOI21 U101 ( .IN1(n74), .IN2(n75), .IN3(n76), .OUT(n77) );
  AOI21 U102 ( .IN1(n821), .IN2(Datain2[8]), .IN3(n77), .OUT(n78) );
  NAND2X1 U103 ( .IN1(n72), .IN2(n78), .OUT(n1095) );
  INVX1 U104 ( .IN(n815), .OUT(n79) );
  NOR2X1 U105 ( .IN1(n1132), .IN2(n79), .OUT(n80) );
  MUX2X1 U106 ( .IN1(add_x_35_A_8_), .IN2(n224), .S(n80), .OUT(n81) );
  NOR2X1 U107 ( .IN1(n1130), .IN2(n81), .OUT(n121) );
  OAI21 U108 ( .IN1(n973), .IN2(add_x_35_A_4_), .IN3(n972), .OUT(n82) );
  NOR2X1 U109 ( .IN1(n957), .IN2(n82), .OUT(n83) );
  AOI22 U110 ( .IN1(n980), .IN2(N159), .IN3(n1034), .IN4(n981), .OUT(n84) );
  NAND2X1 U111 ( .IN1(n83), .IN2(n84), .OUT(n1079) );
  NAND3X1 U112 ( .IN1(n366), .IN2(n382), .IN3(n490), .OUT(n754) );
  INVX1 U113 ( .IN(N159), .OUT(n85) );
  AOI22 U114 ( .IN1(N159), .IN2(DP_OP_982J1_125_6202_n91), .IN3(Datain1[10]), 
        .IN4(n85), .OUT(n86) );
  AOI22 U115 ( .IN1(N159), .IN2(Datain1[9]), .IN3(Datain1[8]), .IN4(n85), 
        .OUT(n87) );
  INVX1 U116 ( .IN(N160), .OUT(n88) );
  AOI22 U117 ( .IN1(N160), .IN2(n86), .IN3(n87), .IN4(n88), .OUT(n89) );
  AOI22 U118 ( .IN1(N159), .IN2(Datain1[15]), .IN3(Datain1[14]), .IN4(n85), 
        .OUT(n90) );
  AOI22 U119 ( .IN1(N159), .IN2(Datain1[13]), .IN3(Datain1[12]), .IN4(n85), 
        .OUT(n91) );
  AOI22 U120 ( .IN1(N160), .IN2(n90), .IN3(n91), .IN4(n88), .OUT(n92) );
  MUX2X1 U121 ( .IN1(n89), .IN2(n92), .S(N161), .OUT(n1189) );
  INVX1 U122 ( .IN(n699), .OUT(n93) );
  INVX1 U123 ( .IN(n698), .OUT(n94) );
  NAND3X1 U124 ( .IN1(n710), .IN2(n93), .IN3(n94), .OUT(n95) );
  INVX1 U125 ( .IN(n719), .OUT(n96) );
  NAND3X1 U126 ( .IN1(n836), .IN2(n95), .IN3(n96), .OUT(n97) );
  INVX1 U127 ( .IN(n713), .OUT(n98) );
  AOI21 U128 ( .IN1(n242), .IN2(n97), .IN3(n98), .OUT(n819) );
  AOI22 U129 ( .IN1(Final_Exponent_reg[0]), .IN2(n647), .IN3(n822), .IN4(
        Datain1[7]), .OUT(n99) );
  INVX1 U130 ( .IN(DP_OP_986_157_3518_n76), .OUT(n100) );
  NAND2X1 U131 ( .IN1(DP_OP_986_157_3518_n50), .IN2(DP_OP_986_157_3518_n56), 
        .OUT(n101) );
  OAI21 U132 ( .IN1(n100), .IN2(n101), .IN3(n650), .OUT(n102) );
  AOI21 U133 ( .IN1(n100), .IN2(n101), .IN3(n102), .OUT(n104) );
  AOI21 U134 ( .IN1(n821), .IN2(Datain2[7]), .IN3(n104), .OUT(n105) );
  NAND2X1 U135 ( .IN1(n99), .IN2(n105), .OUT(n1094) );
  INVX1 U136 ( .IN(n467), .OUT(n106) );
  AOI22 U137 ( .IN1(n537), .IN2(Final_Mantissa_reg[10]), .IN3(Adder_dataout[6]), .IN4(n826), .OUT(n107) );
  OAI21 U138 ( .IN1(n471), .IN2(n545), .IN3(n107), .OUT(n108) );
  AOI21 U139 ( .IN1(n472), .IN2(n491), .IN3(n108), .OUT(n114) );
  INVX1 U140 ( .IN(n232), .OUT(n115) );
  AOI22 U141 ( .IN1(n477), .IN2(n476), .IN3(n478), .IN4(n115), .OUT(n125) );
  AOI22 U142 ( .IN1(n280), .IN2(n473), .IN3(n279), .IN4(n474), .OUT(n126) );
  OAI21 U143 ( .IN1(n209), .IN2(n475), .IN3(n126), .OUT(n127) );
  NAND2X1 U144 ( .IN1(n527), .IN2(n127), .OUT(n128) );
  NAND3X1 U145 ( .IN1(n114), .IN2(n125), .IN3(n128), .OUT(n129) );
  NOR2X1 U146 ( .IN1(n535), .IN2(n536), .OUT(n130) );
  AOI21 U147 ( .IN1(n130), .IN2(n232), .IN3(n129), .OUT(n131) );
  OAI21 U148 ( .IN1(n558), .IN2(n106), .IN3(n131), .OUT(n132) );
  NOR2X1 U149 ( .IN1(n847), .IN2(n551), .OUT(n133) );
  AOI21 U150 ( .IN1(n133), .IN2(n493), .IN3(n132), .OUT(n134) );
  AOI22 U151 ( .IN1(n483), .IN2(n484), .IN3(n485), .IN4(n486), .OUT(n135) );
  AOI22 U152 ( .IN1(n479), .IN2(n480), .IN3(n481), .IN4(n482), .OUT(n136) );
  NAND2X1 U153 ( .IN1(n135), .IN2(n136), .OUT(n137) );
  AOI22 U154 ( .IN1(Final_Mantissa_reg[9]), .IN2(n561), .IN3(n487), .IN4(n137), 
        .OUT(n138) );
  OAI21 U155 ( .IN1(RSTn_BAR), .IN2(n134), .IN3(n138), .OUT(n1063) );
  NAND2X1 U156 ( .IN1(n815), .IN2(n816), .OUT(n139) );
  MUX2X1 U157 ( .IN1(Op2_Mantissa_reg_7_), .IN2(n244), .S(n139), .OUT(n140) );
  NOR2X1 U158 ( .IN1(n1130), .IN2(n140), .OUT(n123) );
  NANDX2 U159 ( .IN1(n722), .IN2(n646), .OUT(C2_Z_0) );
  INVX4 U160 ( .IN(DP_OP_982J1_125_6202_n72), .OUT(N155) );
  NANDX2 U161 ( .IN1(n652), .IN2(n651), .OUT(n1102) );
  NANDX2 U162 ( .IN1(n650), .IN2(C405_DATA2_7), .OUT(n651) );
  INVX1 U163 ( .IN(n562), .OUT(n1062) );
  NAND2X1 U164 ( .IN1(n391), .IN2(n390), .OUT(n1068) );
  NAND2X1 U165 ( .IN1(n819), .IN2(n725), .OUT(n837) );
  NAND2X1 U166 ( .IN1(n528), .IN2(n554), .OUT(n529) );
  NAND2X1 U167 ( .IN1(n494), .IN2(n493), .OUT(n495) );
  INVX1 U168 ( .IN(DP_OP_986_157_3518_n42), .OUT(DP_OP_986_157_3518_n40) );
  NAND2X1 U169 ( .IN1(n419), .IN2(n418), .OUT(n420) );
  NAND2X1 U170 ( .IN1(n441), .IN2(n440), .OUT(n442) );
  INVX1 U171 ( .IN(n724), .OUT(n109) );
  INVX1 U172 ( .IN(n1141), .OUT(n111) );
  NAND2X1 U173 ( .IN1(n824), .IN2(n375), .OUT(n376) );
  NANDX2 U174 ( .IN1(n555), .IN2(n721), .OUT(n383) );
  INVX1 U175 ( .IN(n1143), .OUT(n110) );
  NAND2X1 U176 ( .IN1(n1050), .IN2(n1049), .OUT(n1074) );
  NAND2X1 U177 ( .IN1(n1033), .IN2(n1032), .OUT(n1076) );
  NAND2X1 U178 ( .IN1(n1040), .IN2(n1039), .OUT(n1075) );
  NAND2X1 U179 ( .IN1(n527), .IN2(n408), .OUT(n411) );
  NAND2X1 U180 ( .IN1(n477), .IN2(n409), .OUT(n410) );
  NAND2X1 U181 ( .IN1(n428), .IN2(n427), .OUT(n429) );
  INVX1 U182 ( .IN(n648), .OUT(n649) );
  NANDX2 U183 ( .IN1(n913), .IN2(n912), .OUT(n914) );
  NAND2X1 U184 ( .IN1(n547), .IN2(n546), .OUT(n549) );
  NAND2X1 U185 ( .IN1(n767), .IN2(n766), .OUT(n768) );
  INVX1 U186 ( .IN(n818), .OUT(n124) );
  NANDX2 U187 ( .IN1(n930), .IN2(n929), .OUT(n931) );
  INVX1 U188 ( .IN(n636), .OUT(n661) );
  INVX1 U189 ( .IN(n676), .OUT(n624) );
  INVX1 U190 ( .IN(n1035), .OUT(n1036) );
  INVX1 U191 ( .IN(n1029), .OUT(n1030) );
  NAND2X1 U192 ( .IN1(n769), .IN2(n718), .OUT(n318) );
  NAND2X1 U193 ( .IN1(n492), .IN2(n804), .OUT(n399) );
  INVX1 U194 ( .IN(n804), .OUT(n745) );
  INVX1 U195 ( .IN(n594), .OUT(n761) );
  NANDX2 U196 ( .IN1(n149), .IN2(n150), .OUT(n1167) );
  INVX1 U197 ( .IN(n696), .OUT(n697) );
  INVX1 U198 ( .IN(n669), .OUT(n598) );
  NANDX2 U199 ( .IN1(n146), .IN2(n147), .OUT(n1153) );
  NAND2X1 U200 ( .IN1(n997), .IN2(n996), .OUT(n1003) );
  INVX1 U201 ( .IN(n1129), .OUT(n816) );
  NANDX2 U202 ( .IN1(n1164), .IN2(n151), .OUT(n150) );
  NAND2X1 U203 ( .IN1(n823), .IN2(n578), .OUT(n580) );
  NANDX2 U204 ( .IN1(n1178), .IN2(n154), .OUT(n153) );
  INVX1 U205 ( .IN(n351), .OUT(n267) );
  INVX1 U206 ( .IN(n965), .OUT(n966) );
  INVX1 U207 ( .IN(n1109), .OUT(n1110) );
  NANDX2 U208 ( .IN1(n707), .IN2(n646), .OUT(n696) );
  INVX1 U209 ( .IN(n739), .OUT(n741) );
  NANDX2 U210 ( .IN1(n1150), .IN2(n148), .OUT(n147) );
  INVX1 U211 ( .IN(n1046), .OUT(n1047) );
  NAND2X1 U212 ( .IN1(n536), .IN2(n403), .OUT(n405) );
  INVX1 U213 ( .IN(n764), .OUT(n692) );
  NANDX2 U214 ( .IN1(add_x_35_A_8_), .IN2(n1132), .OUT(n1131) );
  INVX1 U215 ( .IN(n694), .OUT(n612) );
  NANDX2 U216 ( .IN1(n235), .IN2(n691), .OUT(n611) );
  INVX1 U217 ( .IN(n993), .OUT(n964) );
  INVX1 U218 ( .IN(n1015), .OUT(n1017) );
  NAND2X1 U219 ( .IN1(N155), .IN2(n1011), .OUT(n1044) );
  INVX1 U220 ( .IN(n289), .OUT(n1103) );
  NAND2X1 U221 ( .IN1(n740), .IN2(n713), .OUT(n578) );
  NAND2X1 U222 ( .IN1(n280), .IN2(n431), .OUT(n430) );
  INVX1 U223 ( .IN(n535), .OUT(n403) );
  NAND2X1 U224 ( .IN1(N148), .IN2(n984), .OUT(n959) );
  INVX1 U225 ( .IN(n960), .OUT(n923) );
  NANDX2 U226 ( .IN1(n815), .IN2(n499), .OUT(n729) );
  NAND2X1 U227 ( .IN1(n285), .IN2(n565), .OUT(n566) );
  NAND2X1 U228 ( .IN1(n270), .IN2(n157), .OUT(n1111) );
  INVX4 U229 ( .IN(n387), .OUT(n513) );
  INVX1 U230 ( .IN(n896), .OUT(n891) );
  INVX1 U231 ( .IN(n307), .OUT(n308) );
  INVX1 U232 ( .IN(n675), .OUT(n677) );
  INVX1 U233 ( .IN(n601), .OUT(n759) );
  INVX1 U234 ( .IN(n757), .OUT(n683) );
  INVX1 U235 ( .IN(n608), .OUT(n673) );
  NANDX2 U236 ( .IN1(n227), .IN2(n371), .OUT(n722) );
  NAND2X1 U237 ( .IN1(n767), .IN2(n740), .OUT(n719) );
  INVX1 U238 ( .IN(n787), .OUT(Dataout[0]) );
  INVX1 U239 ( .IN(n1130), .OUT(n499) );
  INVX1 U240 ( .IN(n788), .OUT(Dataout[1]) );
  INVX1 U241 ( .IN(n789), .OUT(Dataout[2]) );
  INVX1 U242 ( .IN(n790), .OUT(Dataout[3]) );
  NAND2X1 U243 ( .IN1(n898), .IN2(n1130), .OUT(n288) );
  INVX1 U244 ( .IN(n791), .OUT(Dataout[4]) );
  INVX1 U245 ( .IN(n792), .OUT(Dataout[5]) );
  INVX1 U246 ( .IN(n793), .OUT(Dataout[6]) );
  INVX1 U247 ( .IN(n740), .OUT(n733) );
  INVX1 U248 ( .IN(n794), .OUT(Dataout[7]) );
  INVX1 U249 ( .IN(n795), .OUT(Dataout[8]) );
  INVX1 U250 ( .IN(n796), .OUT(Dataout[9]) );
  INVX1 U251 ( .IN(n797), .OUT(Dataout[10]) );
  INVX1 U252 ( .IN(n798), .OUT(Dataout[11]) );
  INVX1 U253 ( .IN(n799), .OUT(Dataout[12]) );
  INVX1 U254 ( .IN(n801), .OUT(Dataout[13]) );
  INVX1 U255 ( .IN(n820), .OUT(n565) );
  INVX1 U256 ( .IN(n843), .OUT(n845) );
  NANDX2 U257 ( .IN1(add_x_35_A_6_), .IN2(n1134), .OUT(n1133) );
  INVX1 U258 ( .IN(n944), .OUT(n945) );
  INVX1 U259 ( .IN(n774), .OUT(ExcCheck_Datain_1_) );
  INVX1 U260 ( .IN(n779), .OUT(ExcCheck_Datain_6_) );
  INVX4 U261 ( .IN(N364), .OUT(n141) );
  INVX1 U262 ( .IN(N420), .OUT(n142) );
  NAND2X1 U263 ( .IN1(n800), .IN2(Final_Exponent_reg[0]), .OUT(n794) );
  INVX1 U264 ( .IN(n776), .OUT(ExcCheck_Datain_3_) );
  INVX1 U265 ( .IN(n778), .OUT(ExcCheck_Datain_5_) );
  INVX1 U266 ( .IN(n777), .OUT(ExcCheck_Datain_4_) );
  NAND2X1 U267 ( .IN1(n800), .IN2(DP_OP_986_157_3518_n93), .OUT(n797) );
  INVX1 U268 ( .IN(n863), .OUT(n864) );
  INVX1 U269 ( .IN(n773), .OUT(ExcCheck_Datain_0_) );
  NANDX2 U270 ( .IN1(Debug_reg[3]), .IN2(n1144), .OUT(n1139) );
  INVX1 U271 ( .IN(n775), .OUT(ExcCheck_Datain_2_) );
  NAND2X1 U272 ( .IN1(n800), .IN2(n281), .OUT(n792) );
  INVX4 U273 ( .IN(n382), .OUT(n525) );
  NAND2X1 U274 ( .IN1(n800), .IN2(n280), .OUT(n791) );
  NAND2X1 U275 ( .IN1(n800), .IN2(Final_Mantissa_reg[9]), .OUT(n793) );
  NAND2X1 U276 ( .IN1(n800), .IN2(n276), .OUT(n788) );
  NAND2X1 U277 ( .IN1(n800), .IN2(n275), .OUT(n787) );
  NAND2X1 U278 ( .IN1(n800), .IN2(n279), .OUT(n790) );
  INVX1 U279 ( .IN(n736), .OUT(n737) );
  NAND2X1 U280 ( .IN1(n279), .IN2(n306), .OUT(n601) );
  NANDX2 U281 ( .IN1(n328), .IN2(n727), .OUT(n742) );
  NAND2X1 U282 ( .IN1(n868), .IN2(n867), .OUT(n869) );
  INVX1 U283 ( .IN(n802), .OUT(Dataout[14]) );
  INVX1 U284 ( .IN(n618), .OUT(n682) );
  NANDX2 U285 ( .IN1(n284), .IN2(n327), .OUT(n380) );
  INVX1 U286 ( .IN(n316), .OUT(n317) );
  NANDX2 U287 ( .IN1(n588), .IN2(n587), .OUT(n589) );
  INVX1 U288 ( .IN(n854), .OUT(Debug[0]) );
  INVX1 U289 ( .IN(n855), .OUT(Debug[1]) );
  INVX1 U290 ( .IN(n856), .OUT(Debug[2]) );
  INVX1 U291 ( .IN(n860), .OUT(Debug[4]) );
  INVX1 U292 ( .IN(n356), .OUT(n314) );
  INVX1 U293 ( .IN(Dataout_valid), .OUT(n862) );
  NAND2X1 U294 ( .IN1(n281), .IN2(n758), .OUT(n618) );
  NAND2X1 U295 ( .IN1(n1145), .IN2(n285), .OUT(n1147) );
  INVX1 U296 ( .IN(n631), .OUT(n686) );
  NANDX2 U297 ( .IN1(Final_Mantissa_reg[10]), .IN2(n328), .OUT(n708) );
  INVX4 U298 ( .IN(Datain2[10]), .OUT(n178) );
  NAND2X1 U299 ( .IN1(n868), .IN2(Data_valid), .OUT(n884) );
  INVX4 U300 ( .IN(Datain2[11]), .OUT(n179) );
  INVX1 U301 ( .IN(n857), .OUT(Debug[3]) );
  INVX1 U302 ( .IN(n715), .OUT(n716) );
  NAND2X1 U303 ( .IN1(n200), .IN2(DP_OP_982J1_125_6202_n101), .OUT(n184) );
  INVX1 U304 ( .IN(DP_OP_982J1_125_6202_n101), .OUT(n180) );
  INVX4 U305 ( .IN(Datain1[12]), .OUT(n199) );
  INVX4 U306 ( .IN(Datain1[10]), .OUT(n196) );
  INVX4 U307 ( .IN(Datain1[9]), .OUT(n195) );
  NAND2X1 U308 ( .IN1(Final_Exponent_reg[0]), .IN2(DP_OP_986_157_3518_n93), 
        .OUT(n593) );
  NAND2X1 U309 ( .IN1(n275), .IN2(n276), .OUT(n394) );
  NAND2X1 U310 ( .IN1(DP_OP_982J1_125_6202_n102), .IN2(n906), .OUT(n202) );
  NANDX2 U311 ( .IN1(add_x_35_A_2_), .IN2(n1128), .OUT(n1137) );
  BUF4X U312 ( .IN(Final_Exponent_reg[5]), .OUT(n145) );
  INVX1 U313 ( .IN(DP_OP_982J1_125_6202_n102), .OUT(n143) );
  INVX4 U314 ( .IN(DP_OP_982J1_125_6202_n100), .OUT(n144) );
  INVX1 U315 ( .IN(N145), .OUT(n148) );
  NAND2X1 U316 ( .IN1(N145), .IN2(n1151), .OUT(n146) );
  INVX1 U317 ( .IN(N149), .OUT(n151) );
  NAND2X1 U318 ( .IN1(N149), .IN2(n1165), .OUT(n149) );
  NAND2X1 U319 ( .IN1(n152), .IN2(n153), .OUT(n1181) );
  INVX1 U320 ( .IN(N153), .OUT(n154) );
  NAND2X1 U321 ( .IN1(N153), .IN2(n1179), .OUT(n152) );
  INVX4 U322 ( .IN(n155), .OUT(n156) );
  INVX4 U323 ( .IN(N143), .OUT(n157) );
  NAND2X1 U324 ( .IN1(DP_OP_986_157_3518_n38), .IN2(n158), .OUT(
        DP_OP_986_157_3518_n12) );
  NAND2X1 U325 ( .IN1(DP_OP_986_157_3518_n28), .IN2(n159), .OUT(
        DP_OP_986_157_3518_n2) );
  NAND2X1 U326 ( .IN1(C1_Z_3), .IN2(n160), .OUT(DP_OP_986_157_3518_n62) );
  NAND2X1 U327 ( .IN1(C1_Z_2), .IN2(n161), .OUT(DP_OP_986_157_3518_n66) );
  INVX1 U328 ( .IN(DP_OP_986_157_3518_n36), .OUT(DP_OP_986_157_3518_n53) );
  NANDX2 U329 ( .IN1(n166), .IN2(DP_OP_986_157_3518_n70), .OUT(
        DP_OP_986_157_3518_n72) );
  NANDX2 U330 ( .IN1(DP_OP_986_157_3518_n50), .IN2(n164), .OUT(n165) );
  NANDX2 U331 ( .IN1(n165), .IN2(n168), .OUT(n169) );
  NANDX2 U332 ( .IN1(DP_OP_986_157_3518_n45), .IN2(n169), .OUT(
        DP_OP_986_157_3518_n43) );
  INVX4 U333 ( .IN(DP_OP_986_157_3518_n33), .OUT(DP_OP_986_157_3518_n52) );
  INVX4 U334 ( .IN(DP_OP_986_157_3518_n30), .OUT(DP_OP_986_157_3518_n51) );
  NANDX2 U335 ( .IN1(DP_OP_986_157_3518_n7), .IN2(DP_OP_986_157_3518_n28), 
        .OUT(n159) );
  NANDX2 U336 ( .IN1(DP_OP_986_157_3518_n7), .IN2(n159), .OUT(
        DP_OP_986_157_3518_n1) );
  NANDX2 U337 ( .IN1(C2_Z_0), .IN2(C1_Z_3), .OUT(n160) );
  NANDX2 U338 ( .IN1(C2_Z_0), .IN2(n160), .OUT(DP_OP_986_157_3518_n61) );
  NANDX2 U339 ( .IN1(n239), .IN2(n167), .OUT(n168) );
  NANDX2 U340 ( .IN1(C2_Z_0), .IN2(C1_Z_2), .OUT(n161) );
  NANDX2 U341 ( .IN1(C2_Z_0), .IN2(C1_Z_1), .OUT(n162) );
  NANDX2 U342 ( .IN1(C2_Z_0), .IN2(C1_Z_0), .OUT(n163) );
  NANDX2 U343 ( .IN1(C2_Z_0), .IN2(n162), .OUT(n166) );
  NANDX2 U344 ( .IN1(DP_OP_986_157_3518_n56), .IN2(DP_OP_986_157_3518_n76), 
        .OUT(n164) );
  NANDX2 U345 ( .IN1(C2_Z_0), .IN2(n161), .OUT(DP_OP_986_157_3518_n65) );
  NAND2X1 U346 ( .IN1(DP_OP_986_157_3518_n24), .IN2(DP_OP_986_157_3518_n38), 
        .OUT(n158) );
  INVX1 U347 ( .IN(DP_OP_986_157_3518_n34), .OUT(DP_OP_986_157_3518_n32) );
  INVX4 U348 ( .IN(DP_OP_986_157_3518_n49), .OUT(DP_OP_986_157_3518_n56) );
  INVX4 U349 ( .IN(DP_OP_986_157_3518_n72), .OUT(n167) );
  NANDX2 U350 ( .IN1(C1_Z_1), .IN2(n162), .OUT(DP_OP_986_157_3518_n70) );
  INVX1 U351 ( .IN(DP_OP_986_157_3518_n41), .OUT(DP_OP_986_157_3518_n54) );
  NAND2X1 U352 ( .IN1(DP_OP_986_157_3518_n24), .IN2(n158), .OUT(
        DP_OP_986_157_3518_n11) );
  MUX2X1 U353 ( .IN1(Datain1[7]), .IN2(n181), .S(Datain2[7]), .OUT(N147) );
  AOI22 U354 ( .IN1(N363), .IN2(N143), .IN3(N147), .IN4(N148), .OUT(N144) );
  NOR2X1 U355 ( .IN1(N148), .IN2(N143), .OUT(n170) );
  MUX2X1 U356 ( .IN1(n141), .IN2(N364), .S(n170), .OUT(N153) );
  AOI21 U357 ( .IN1(n157), .IN2(N363), .IN3(N364), .OUT(n171) );
  MUX2X1 U358 ( .IN1(N365), .IN2(n182), .S(n171), .OUT(N154) );
  AOI22 U359 ( .IN1(N364), .IN2(N148), .IN3(N363), .IN4(n141), .OUT(N149) );
  MUX2X1 U360 ( .IN1(n182), .IN2(N365), .S(n172), .OUT(N150) );
  NOR2X1 U361 ( .IN1(N363), .IN2(N147), .OUT(n173) );
  MUX2X1 U362 ( .IN1(N364), .IN2(n141), .S(n173), .OUT(N145) );
  NAND3X1 U363 ( .IN1(N148), .IN2(N143), .IN3(n141), .OUT(n174) );
  MUX2X1 U364 ( .IN1(n182), .IN2(N365), .S(n174), .OUT(N146) );
  MUX2X1 U365 ( .IN1(DP_OP_982J1_125_6202_n102), .IN2(n143), .S(
        DP_OP_981J1_124_6202_n49), .OUT(n175) );
  MUX2X1 U366 ( .IN1(n906), .IN2(Datain1[14]), .S(n175), .OUT(N369) );
  MUX2X1 U367 ( .IN1(DP_OP_982J1_125_6202_n101), .IN2(n180), .S(n200), .OUT(
        n187) );
  MUX2X1 U368 ( .IN1(DP_OP_981J1_124_6202_n50), .IN2(n186), .S(n187), .OUT(
        N368) );
  INVX1 U369 ( .IN(N365), .OUT(n182) );
  INVX1 U370 ( .IN(DP_OP_981J1_124_6202_n50), .OUT(n186) );
  NAND2X1 U371 ( .IN1(Datain1[13]), .IN2(n180), .OUT(n183) );
  INVX4 U372 ( .IN(Datain1[7]), .OUT(n181) );
  INVX4 U373 ( .IN(Datain2[8]), .OUT(n176) );
  NANDX2 U374 ( .IN1(Datain2[7]), .IN2(n181), .OUT(DP_OP_981J1_124_6202_n55)
         );
  INVX4 U375 ( .IN(DP_OP_982J1_125_6202_n97), .OUT(n177) );
  NANDX2 U376 ( .IN1(n183), .IN2(n185), .OUT(DP_OP_981J1_124_6202_n49) );
  INVX4 U377 ( .IN(N147), .OUT(N143) );
  INVX4 U378 ( .IN(N144), .OUT(N152) );
  NANDX2 U379 ( .IN1(n184), .IN2(DP_OP_981J1_124_6202_n50), .OUT(n185) );
  INVX4 U380 ( .IN(N363), .OUT(N148) );
  NANDX2 U381 ( .IN1(N148), .IN2(n141), .OUT(n172) );
  MUX2X1 U382 ( .IN1(Datain2[7]), .IN2(n193), .S(Datain1[7]), .OUT(
        DP_OP_982J1_125_6202_n72) );
  AOI22 U383 ( .IN1(N419), .IN2(N155), .IN3(N159), .IN4(N160), .OUT(N156) );
  NOR2X1 U384 ( .IN1(N160), .IN2(N155), .OUT(n188) );
  MUX2X1 U385 ( .IN1(n142), .IN2(N420), .S(n188), .OUT(N165) );
  AOI21 U386 ( .IN1(N159), .IN2(N419), .IN3(N420), .OUT(n189) );
  MUX2X1 U387 ( .IN1(N421), .IN2(n197), .S(n189), .OUT(N166) );
  AOI22 U388 ( .IN1(N420), .IN2(N160), .IN3(N419), .IN4(n142), .OUT(N161) );
  NAND2X1 U389 ( .IN1(N160), .IN2(n142), .OUT(n190) );
  MUX2X1 U390 ( .IN1(n197), .IN2(N421), .S(n190), .OUT(N162) );
  NOR2X1 U391 ( .IN1(N419), .IN2(N159), .OUT(n191) );
  MUX2X1 U392 ( .IN1(N420), .IN2(n142), .S(n191), .OUT(N157) );
  NAND3X1 U393 ( .IN1(N160), .IN2(N155), .IN3(n142), .OUT(n192) );
  MUX2X1 U394 ( .IN1(n197), .IN2(N421), .S(n192), .OUT(N158) );
  MUX2X1 U395 ( .IN1(n143), .IN2(DP_OP_982J1_125_6202_n102), .S(Datain1[14]), 
        .OUT(n201) );
  OAI21 U396 ( .IN1(DP_OP_982J1_125_6202_n102), .IN2(n906), .IN3(n202), .OUT(
        n203) );
  MUX2X1 U397 ( .IN1(n201), .IN2(n203), .S(DP_OP_982J1_125_6202_n49), .OUT(
        N425) );
  INVX1 U398 ( .IN(N421), .OUT(n197) );
  INVX1 U399 ( .IN(Datain1[13]), .OUT(n200) );
  INVX4 U400 ( .IN(Datain2[7]), .OUT(n193) );
  INVX4 U401 ( .IN(Datain1[8]), .OUT(n194) );
  NANDX2 U402 ( .IN1(Datain1[7]), .IN2(n193), .OUT(DP_OP_982J1_125_6202_n55)
         );
  INVX4 U403 ( .IN(DP_OP_982J1_125_6202_n91), .OUT(n198) );
  INVX4 U404 ( .IN(N156), .OUT(N164) );
  INVX4 U405 ( .IN(N155), .OUT(N159) );
  INVX4 U406 ( .IN(N419), .OUT(N160) );
  NAND2X1 U407 ( .IN1(n370), .IN2(n657), .OUT(n466) );
  NAND2X1 U408 ( .IN1(n235), .IN2(n674), .OUT(n620) );
  NAND2X1 U409 ( .IN1(n650), .IN2(C405_DATA2_3), .OUT(n584) );
  INVX4 U410 ( .IN(n602), .OUT(n752) );
  NAND2X1 U411 ( .IN1(carry_reg), .IN2(n371), .OUT(n762) );
  NANDX2 U412 ( .IN1(n727), .IN2(n751), .OUT(n767) );
  NANDX2 U413 ( .IN1(n508), .IN2(n507), .OUT(n113) );
  INVX4 U414 ( .IN(n1118), .OUT(n821) );
  NANDX2 U415 ( .IN1(n827), .IN2(n564), .OUT(n535) );
  NANDX2 U416 ( .IN1(n271), .IN2(n1038), .OUT(n269) );
  NANDX2 U417 ( .IN1(n280), .IN2(n758), .OUT(n316) );
  NAND2X1 U418 ( .IN1(n283), .IN2(n313), .OUT(n594) );
  BUF4X U419 ( .IN(Final_Mantissa_reg[1]), .OUT(n283) );
  INVX1 U420 ( .IN(n754), .OUT(n656) );
  INVX1 U421 ( .IN(n998), .OUT(n1120) );
  INVX1 U422 ( .IN(n617), .OUT(n630) );
  INVX4 U423 ( .IN(n1116), .OUT(n822) );
  INVX4 U424 ( .IN(n755), .OUT(n665) );
  NANDX2 U425 ( .IN1(n349), .IN2(n348), .OUT(n755) );
  NANDX2 U426 ( .IN1(n471), .IN2(n544), .OUT(n556) );
  NANDX2 U427 ( .IN1(n267), .IN2(n348), .OUT(n266) );
  NAND2X1 U428 ( .IN1(n209), .IN2(n231), .OUT(n253) );
  NAND2X1 U429 ( .IN1(n278), .IN2(n452), .OUT(n451) );
  NAND2X1 U430 ( .IN1(n485), .IN2(n749), .OUT(n662) );
  INVX4 U431 ( .IN(n266), .OUT(n659) );
  NAND2X1 U432 ( .IN1(n282), .IN2(n238), .OUT(n356) );
  NANDX2 U433 ( .IN1(n210), .IN2(n334), .OUT(n327) );
  BUF8X U434 ( .IN(Final_Mantissa_reg[2]), .OUT(n284) );
  INVX1 U435 ( .IN(Datain1[14]), .OUT(n906) );
  NANDX2 U436 ( .IN1(n490), .IN2(n486), .OUT(n393) );
  NANDX2 U437 ( .IN1(n546), .IN2(n527), .OUT(n502) );
  NAND2X1 U438 ( .IN1(n272), .IN2(Exc_Ack), .OUT(n835) );
  NANDX2 U439 ( .IN1(n822), .IN2(n1112), .OUT(n985) );
  INVX4 U440 ( .IN(n621), .OUT(n658) );
  INVX4 U441 ( .IN(n556), .OUT(n749) );
  INVX4 U442 ( .IN(n327), .OUT(n326) );
  NANDX2 U443 ( .IN1(n481), .IN2(n544), .OUT(n256) );
  NANDX2 U444 ( .IN1(n206), .IN2(n262), .OUT(n259) );
  NAND2X1 U445 ( .IN1(n869), .IN2(n220), .OUT(n870) );
  NAND2X1 U446 ( .IN1(n282), .IN2(n506), .OUT(n507) );
  NANDX2 U447 ( .IN1(n718), .IN2(n320), .OUT(n475) );
  NANDX2 U448 ( .IN1(n769), .IN2(n321), .OUT(n319) );
  NANDX2 U449 ( .IN1(n385), .IN2(n384), .OUT(n386) );
  INVX4 U450 ( .IN(n1138), .OUT(n826) );
  NANDX2 U451 ( .IN1(n273), .IN2(N155), .OUT(n965) );
  NANDX2 U452 ( .IN1(n978), .IN2(n822), .OUT(n924) );
  BUF4X U453 ( .IN(n866), .OUT(n272) );
  NANDX2 U454 ( .IN1(n686), .IN2(n660), .OUT(n632) );
  NANDX2 U455 ( .IN1(n235), .IN2(n681), .OUT(n660) );
  INVX4 U456 ( .IN(n365), .OUT(n367) );
  NANDX2 U457 ( .IN1(n208), .IN2(n326), .OUT(n345) );
  INVX4 U458 ( .IN(n253), .OUT(n252) );
  INVX4 U459 ( .IN(n256), .OUT(n255) );
  NANDX2 U460 ( .IN1(n205), .IN2(n338), .OUT(n353) );
  NANDX2 U461 ( .IN1(n337), .IN2(n341), .OUT(n338) );
  INVX4 U462 ( .IN(n340), .OUT(n341) );
  NANDX2 U463 ( .IN1(n231), .IN2(n254), .OUT(n340) );
  INVX4 U464 ( .IN(n259), .OUT(n258) );
  NANDX2 U465 ( .IN1(n336), .IN2(n261), .OUT(n257) );
  NANDX2 U466 ( .IN1(n233), .IN2(n210), .OUT(n263) );
  NANDX2 U467 ( .IN1(n815), .IN2(n708), .OUT(n298) );
  INVX4 U468 ( .IN(n582), .OUT(n577) );
  INVX4 U469 ( .IN(RSTn_BAR), .OUT(n285) );
  INVX4 U470 ( .IN(n786), .OUT(ExcCheck_Datain_14_) );
  INVX4 U471 ( .IN(n785), .OUT(ExcCheck_Datain_12_) );
  INVX4 U472 ( .IN(n784), .OUT(ExcCheck_Datain_11_) );
  INVX4 U473 ( .IN(n782), .OUT(ExcCheck_Datain_9_) );
  INVX4 U474 ( .IN(n781), .OUT(ExcCheck_Datain_8_) );
  INVX1 U475 ( .IN(Datain2[15]), .OUT(n293) );
  INVX1 U476 ( .IN(Datain1[15]), .OUT(n295) );
  NANDX2 U477 ( .IN1(n717), .IN2(n716), .OUT(n1144) );
  INVX4 U478 ( .IN(n510), .OUT(n515) );
  INVX4 U479 ( .IN(n509), .OUT(n521) );
  NANDX2 U480 ( .IN1(n527), .IN2(n548), .OUT(n530) );
  NANDX2 U481 ( .IN1(n426), .IN2(n425), .OUT(n510) );
  NANDX2 U482 ( .IN1(n424), .IN2(n423), .OUT(n509) );
  NANDX2 U483 ( .IN1(n393), .IN2(n392), .OUT(n528) );
  NANDX2 U484 ( .IN1(n389), .IN2(n388), .OUT(n417) );
  INVX4 U485 ( .IN(n558), .OUT(n439) );
  INVX4 U486 ( .IN(n409), .OUT(n333) );
  NANDX2 U487 ( .IN1(n324), .IN2(n323), .OUT(n409) );
  INVX4 U488 ( .IN(n520), .OUT(n487) );
  NANDX2 U489 ( .IN1(n285), .IN2(n554), .OUT(n520) );
  NANDX2 U490 ( .IN1(n449), .IN2(n448), .OUT(n476) );
  INVX4 U491 ( .IN(n459), .OUT(n477) );
  NANDX2 U492 ( .IN1(n739), .IN2(n492), .OUT(n459) );
  INVX4 U493 ( .IN(n318), .OUT(n474) );
  INVX4 U494 ( .IN(n516), .OUT(n527) );
  NANDX2 U495 ( .IN1(n492), .IN2(n315), .OUT(n516) );
  INVX4 U496 ( .IN(n399), .OUT(n472) );
  NANDX2 U497 ( .IN1(n447), .IN2(n446), .OUT(n467) );
  INVX4 U498 ( .IN(n383), .OUT(n479) );
  INVX4 U499 ( .IN(n381), .OUT(n482) );
  NANDX2 U500 ( .IN1(n466), .IN2(n494), .OUT(n558) );
  NANDX2 U501 ( .IN1(n397), .IN2(n396), .OUT(n548) );
  INVX4 U502 ( .IN(n475), .OUT(n450) );
  INVX4 U503 ( .IN(n319), .OUT(n473) );
  INVX4 U504 ( .IN(n322), .OUT(n546) );
  NANDX2 U505 ( .IN1(n321), .IN2(n320), .OUT(n322) );
  INVX4 U506 ( .IN(n769), .OUT(n320) );
  INVX4 U507 ( .IN(n718), .OUT(n321) );
  INVX4 U508 ( .IN(n523), .OUT(n537) );
  INVX4 U509 ( .IN(n567), .OUT(n561) );
  NANDX2 U510 ( .IN1(n721), .IN2(n384), .OUT(n505) );
  INVX4 U511 ( .IN(n385), .OUT(n721) );
  INVX4 U512 ( .IN(n386), .OUT(n486) );
  INVX4 U513 ( .IN(n555), .OUT(n384) );
  NANDX2 U514 ( .IN1(n657), .IN2(n369), .OUT(n555) );
  NANDX2 U515 ( .IN1(n657), .IN2(n364), .OUT(n385) );
  INVX4 U516 ( .IN(n376), .OUT(n494) );
  INVX4 U517 ( .IN(n747), .OUT(n375) );
  NANDX2 U518 ( .IN1(n750), .IN2(n400), .OUT(n747) );
  INVX4 U519 ( .IN(n470), .OUT(n491) );
  NANDX2 U520 ( .IN1(n469), .IN2(n468), .OUT(n470) );
  NANDX2 U521 ( .IN1(n694), .IN2(n308), .OUT(n739) );
  INVX4 U522 ( .IN(n437), .OUT(n492) );
  INVX4 U523 ( .IN(n545), .OUT(n526) );
  NANDX2 U524 ( .IN1(n717), .IN2(n567), .OUT(n533) );
  NANDX2 U525 ( .IN1(n897), .IN2(n715), .OUT(n567) );
  NANDX2 U526 ( .IN1(n285), .IN2(n827), .OUT(n717) );
  INVX4 U527 ( .IN(n670), .OUT(n710) );
  NANDX2 U528 ( .IN1(n686), .IN2(n685), .OUT(n687) );
  INVX4 U529 ( .IN(n680), .OUT(n689) );
  NANDX2 U530 ( .IN1(n679), .IN2(n678), .OUT(n680) );
  NANDX2 U531 ( .IN1(n677), .IN2(n676), .OUT(n678) );
  NANDX2 U532 ( .IN1(n668), .IN2(n667), .OUT(n836) );
  INVX4 U533 ( .IN(n706), .OUT(n667) );
  INVX4 U534 ( .IN(n660), .OUT(n685) );
  INVX4 U535 ( .IN(n655), .OUT(n690) );
  NANDX2 U536 ( .IN1(n564), .IN2(n563), .OUT(n1125) );
  INVX4 U537 ( .IN(n402), .OUT(n431) );
  NANDX2 U538 ( .IN1(n279), .IN2(n395), .OUT(n402) );
  INVX4 U539 ( .IN(n451), .OUT(n395) );
  INVX4 U540 ( .IN(n394), .OUT(n452) );
  INVX4 U541 ( .IN(n380), .OUT(n564) );
  NAND2X1 U542 ( .IN1(Datain2[10]), .IN2(n821), .OUT(n585) );
  NANDX2 U543 ( .IN1(n500), .IN2(n1115), .OUT(n1071) );
  INVX4 U544 ( .IN(n1052), .OUT(n973) );
  INVX4 U545 ( .IN(n958), .OUT(n981) );
  INVX4 U546 ( .IN(n1020), .OUT(n1022) );
  INVX4 U547 ( .IN(n729), .OUT(n817) );
  NANDX2 U548 ( .IN1(n947), .IN2(n946), .OUT(n948) );
  INVX4 U549 ( .IN(n1055), .OUT(n1045) );
  NANDX2 U550 ( .IN1(N160), .IN2(n1038), .OUT(n1055) );
  INVX4 U551 ( .IN(n269), .OUT(n1019) );
  INVX4 U552 ( .IN(n924), .OUT(n1053) );
  NANDX2 U553 ( .IN1(n1146), .IN2(n579), .OUT(n1052) );
  NANDX2 U554 ( .IN1(n917), .IN2(n942), .OUT(n1031) );
  INVX1 U555 ( .IN(Datain1[6]), .OUT(n1011) );
  NANDX2 U556 ( .IN1(n821), .IN2(n944), .OUT(n1001) );
  NANDX2 U557 ( .IN1(n910), .IN2(n909), .OUT(n944) );
  INVX4 U558 ( .IN(n287), .OUT(n825) );
  NAND2X1 U559 ( .IN1(n286), .IN2(n204), .OUT(n287) );
  NAND2X1 U560 ( .IN1(StateMC[0]), .IN2(StateMC[1]), .OUT(n851) );
  NAND2X1 U561 ( .IN1(StateMC[0]), .IN2(StateMC[2]), .OUT(n1058) );
  NAND2X1 U562 ( .IN1(StateMC[1]), .IN2(n204), .OUT(n897) );
  NANDX2 U563 ( .IN1(n142), .IN2(n999), .OUT(n998) );
  INVX4 U564 ( .IN(n1051), .OUT(n1117) );
  NANDX2 U565 ( .IN1(n1112), .IN2(N148), .OUT(n1051) );
  NANDX2 U566 ( .IN1(n141), .IN2(n932), .OUT(n268) );
  NANDX2 U567 ( .IN1(n303), .IN2(n306), .OUT(n757) );
  INVX4 U568 ( .IN(n632), .OUT(n634) );
  INVX4 U569 ( .IN(n663), .OUT(n681) );
  NANDX2 U570 ( .IN1(n630), .IN2(n629), .OUT(C1_Z_1) );
  NANDX2 U571 ( .IN1(n355), .IN2(n662), .OUT(n621) );
  NANDX2 U572 ( .IN1(n620), .IN2(n663), .OUT(n676) );
  INVX4 U573 ( .IN(n607), .OUT(n674) );
  NANDX2 U574 ( .IN1(n695), .IN2(n614), .OUT(n643) );
  NANDX2 U575 ( .IN1(n275), .IN2(n310), .OUT(n694) );
  NANDX2 U576 ( .IN1(n370), .IN2(n352), .OUT(n657) );
  NANDX2 U577 ( .IN1(n264), .IN2(n348), .OUT(n370) );
  INVX4 U578 ( .IN(n666), .OUT(n695) );
  NANDX2 U579 ( .IN1(n611), .IN2(n610), .OUT(n666) );
  INVX4 U580 ( .IN(n748), .OUT(n348) );
  NANDX2 U581 ( .IN1(n544), .IN2(n362), .OUT(n748) );
  INVX4 U582 ( .IN(n359), .OUT(n445) );
  NANDX2 U583 ( .IN1(n305), .IN2(n306), .OUT(n608) );
  INVX4 U584 ( .IN(n671), .OUT(n610) );
  NANDX2 U585 ( .IN1(n607), .IN2(n606), .OUT(n671) );
  NANDX2 U586 ( .IN1(n239), .IN2(n691), .OUT(n606) );
  NANDX2 U587 ( .IN1(n207), .IN2(n691), .OUT(n607) );
  INVX4 U588 ( .IN(n372), .OUT(n654) );
  NANDX2 U589 ( .IN1(n367), .IN2(n366), .OUT(n372) );
  NANDX2 U590 ( .IN1(n314), .IN2(n313), .OUT(n669) );
  NANDX2 U591 ( .IN1(n655), .IN2(n596), .OUT(n644) );
  INVX4 U592 ( .IN(n312), .OUT(n313) );
  NANDX2 U593 ( .IN1(n311), .IN2(n310), .OUT(n312) );
  INVX4 U594 ( .IN(n373), .OUT(n366) );
  NANDX2 U595 ( .IN1(n357), .IN2(n356), .OUT(n490) );
  NANDX2 U596 ( .IN1(n593), .IN2(n653), .OUT(n655) );
  INVX4 U597 ( .IN(n704), .OUT(n653) );
  NANDX2 U598 ( .IN1(n592), .IN2(n591), .OUT(n704) );
  NANDX2 U599 ( .IN1(n347), .IN2(n346), .OUT(n398) );
  NANDX2 U600 ( .IN1(n335), .IN2(n345), .OUT(n387) );
  NANDX2 U601 ( .IN1(n255), .IN2(n362), .OUT(n602) );
  INVX4 U602 ( .IN(n344), .OUT(n362) );
  NANDX2 U603 ( .IN1(n343), .IN2(n471), .OUT(n344) );
  NANDX2 U604 ( .IN1(n252), .IN2(n254), .OUT(n342) );
  INVX4 U605 ( .IN(n360), .OUT(n544) );
  INVX4 U606 ( .IN(n339), .OUT(n254) );
  NANDX2 U607 ( .IN1(n260), .IN2(n258), .OUT(n339) );
  NANDX2 U608 ( .IN1(n262), .IN2(n260), .OUT(n347) );
  INVX4 U609 ( .IN(n257), .OUT(n260) );
  INVX4 U610 ( .IN(n263), .OUT(n262) );
  BUF4X U611 ( .IN(N691), .OUT(n282) );
  NANDX2 U612 ( .IN1(n309), .IN2(n310), .OUT(n764) );
  INVX4 U613 ( .IN(n302), .OUT(n310) );
  NANDX2 U614 ( .IN1(n301), .IN2(n306), .OUT(n302) );
  INVX4 U615 ( .IN(n738), .OUT(n306) );
  NANDX2 U616 ( .IN1(n300), .IN2(n758), .OUT(n738) );
  INVX4 U617 ( .IN(n299), .OUT(n758) );
  BUF4X U618 ( .IN(Final_Mantissa_reg[3]), .OUT(n275) );
  INVX4 U619 ( .IN(n590), .OUT(n691) );
  NANDX2 U620 ( .IN1(n234), .IN2(n591), .OUT(n590) );
  INVX4 U621 ( .IN(n589), .OUT(n591) );
  INVX4 U622 ( .IN(n805), .OUT(n646) );
  NANDX2 U623 ( .IN1(n742), .IN2(n762), .OUT(n805) );
  NANDX2 U624 ( .IN1(n582), .IN2(n581), .OUT(n707) );
  INVX4 U625 ( .IN(n298), .OUT(n371) );
  NANDX2 U626 ( .IN1(n580), .IN2(n579), .OUT(n647) );
  NANDX2 U627 ( .IN1(n577), .IN2(n581), .OUT(n713) );
  INVX4 U628 ( .IN(n767), .OUT(n581) );
  NANDX2 U629 ( .IN1(n576), .IN2(n575), .OUT(n582) );
  BUF4X U630 ( .IN(Final_Exponent_reg[3]), .OUT(DP_OP_986_157_3518_n93) );
  NANDX2 U631 ( .IN1(n297), .IN2(n296), .OUT(n815) );
  NAND2X1 U632 ( .IN1(Op1_Sign_reg), .IN2(n229), .OUT(n296) );
  NAND2X1 U633 ( .IN1(Op2_Sign_reg), .IN2(n228), .OUT(n297) );
  NANDX2 U634 ( .IN1(n885), .IN2(n291), .OUT(n1118) );
  BUF4X U635 ( .IN(Datain2[9]), .OUT(DP_OP_982J1_125_6202_n97) );
  BUF4X U636 ( .IN(Datain2[12]), .OUT(DP_OP_982J1_125_6202_n100) );
  BUF4X U637 ( .IN(Datain2[13]), .OUT(DP_OP_982J1_125_6202_n101) );
  BUF4X U638 ( .IN(Datain2[14]), .OUT(DP_OP_982J1_125_6202_n102) );
  NAND2X1 U639 ( .IN1(n204), .IN2(n220), .OUT(n846) );
  INVX1 U640 ( .IN(n824), .OUT(n847) );
  NAND2X1 U641 ( .IN1(n815), .IN2(n1137), .OUT(n813) );
  NAND2X1 U642 ( .IN1(n815), .IN2(n1135), .OUT(n811) );
  NAND2X1 U643 ( .IN1(Dataout_valid), .IN2(Final_Exponent_reg[7]), .OUT(n802)
         );
  NAND2X1 U644 ( .IN1(n800), .IN2(n278), .OUT(n789) );
  NAND2X1 U645 ( .IN1(n800), .IN2(Final_Exponent_reg[4]), .OUT(n798) );
  NAND2X1 U646 ( .IN1(n800), .IN2(Final_Exponent_reg[2]), .OUT(n796) );
  NAND2X1 U647 ( .IN1(n800), .IN2(Final_Exponent_reg[1]), .OUT(n795) );
  NAND2X1 U648 ( .IN1(n800), .IN2(n145), .OUT(n799) );
  NAND2X1 U649 ( .IN1(n800), .IN2(n156), .OUT(n801) );
  NAND2X1 U650 ( .IN1(n815), .IN2(n1133), .OUT(n809) );
  NAND2X1 U651 ( .IN1(n735), .IN2(n824), .OUT(n736) );
  NAND2X1 U652 ( .IN1(n815), .IN2(n762), .OUT(n734) );
  NAND2X1 U653 ( .IN1(n815), .IN2(n1131), .OUT(n807) );
  NAND2X1 U654 ( .IN1(n278), .IN2(n518), .OUT(n463) );
  INVX1 U655 ( .IN(n714), .OUT(n894) );
  INVX1 U656 ( .IN(n398), .OUT(n456) );
  NAND2X1 U657 ( .IN1(n385), .IN2(n555), .OUT(n381) );
  NAND2X1 U658 ( .IN1(n282), .IN2(n473), .OUT(n397) );
  INVX1 U659 ( .IN(n803), .OUT(n551) );
  NAND2X1 U660 ( .IN1(n754), .IN2(n372), .OUT(n374) );
  NAND2X1 U661 ( .IN1(n824), .IN2(n805), .OUT(n437) );
  NAND2X1 U662 ( .IN1(n824), .IN2(n581), .OUT(n523) );
  NAND2X1 U663 ( .IN1(n824), .IN2(n733), .OUT(n545) );
  INVX1 U664 ( .IN(n711), .OUT(n700) );
  NAND2X1 U665 ( .IN1(n708), .IN2(n707), .OUT(n709) );
  NAND2X1 U666 ( .IN1(Final_Mantissa_reg[10]), .IN2(Final_Mantissa_reg[9]), 
        .OUT(n534) );
  INVX1 U667 ( .IN(n851), .OUT(n726) );
  BUF4X U668 ( .IN(N419), .OUT(n271) );
  BUF4X U669 ( .IN(Datain1[5]), .OUT(n273) );
  BUF4X U670 ( .IN(N363), .OUT(n270) );
  INVX4 U671 ( .IN(n268), .OUT(n1112) );
  INVX1 U672 ( .IN(n616), .OUT(C1_Z_2) );
  INVX1 U673 ( .IN(n640), .OUT(n641) );
  NAND2X1 U674 ( .IN1(n353), .IN2(n483), .OUT(n636) );
  INVX1 U675 ( .IN(n471), .OUT(n483) );
  NAND2X1 U676 ( .IN1(Final_Mantissa_reg[9]), .IN2(n205), .OUT(n631) );
  INVX1 U677 ( .IN(n742), .OUT(n635) );
  INVX1 U678 ( .IN(n480), .OUT(n354) );
  NAND2X1 U679 ( .IN1(n209), .IN2(n317), .OUT(n675) );
  INVX1 U680 ( .IN(n662), .OUT(n619) );
  NAND2X1 U681 ( .IN1(n612), .IN2(n805), .OUT(n613) );
  NAND2X1 U682 ( .IN1(n265), .IN2(n351), .OUT(n264) );
  INVX1 U683 ( .IN(n481), .OUT(n350) );
  INVX1 U684 ( .IN(n600), .OUT(C1_Z_3) );
  NAND2X1 U685 ( .IN1(n805), .IN2(n761), .OUT(n595) );
  NAND2X1 U686 ( .IN1(n283), .IN2(n236), .OUT(n357) );
  INVX1 U687 ( .IN(n334), .OUT(n358) );
  NAND2X1 U688 ( .IN1(n205), .IN2(n232), .OUT(n299) );
  NAND2X1 U689 ( .IN1(n206), .IN2(n237), .OUT(n304) );
  INVX1 U690 ( .IN(n328), .OUT(n751) );
  NAND2X1 U691 ( .IN1(Final_Exponent_reg[4]), .IN2(Final_Exponent_reg[7]), 
        .OUT(n573) );
  NAND2X1 U692 ( .IN1(Final_Exponent_reg[6]), .IN2(n145), .OUT(n574) );
  NAND2X1 U693 ( .IN1(Final_Exponent_reg[2]), .IN2(DP_OP_986_157_3518_n93), 
        .OUT(n571) );
  NAND2X1 U694 ( .IN1(Final_Exponent_reg[0]), .IN2(Final_Exponent_reg[1]), 
        .OUT(n572) );
  NAND2X1 U695 ( .IN1(n815), .IN2(n325), .OUT(n740) );
  INVX1 U696 ( .IN(n708), .OUT(n325) );
  INVX1 U697 ( .IN(n840), .OUT(n290) );
  INVX1 U698 ( .IN(n886), .OUT(n291) );
  BUF4X U699 ( .IN(Datain1[11]), .OUT(DP_OP_982J1_125_6202_n91) );
  BUF4X U700 ( .IN(Final_Mantissa_reg[6]), .OUT(n279) );
  BUF4X U701 ( .IN(Final_Mantissa_reg[8]), .OUT(n281) );
  BUF4X U702 ( .IN(Final_Mantissa_reg[7]), .OUT(n280) );
  BUF4X U703 ( .IN(Final_Mantissa_reg[4]), .OUT(n276) );
  BUF4X U704 ( .IN(Final_Mantissa_reg[5]), .OUT(n278) );
  NOR2X1 U705 ( .IN1(n284), .IN2(n283), .OUT(n261) );
  NOR2X1 U706 ( .IN1(n481), .IN2(n349), .OUT(n265) );
  TIEHI U707 ( .OUT(n73) );
  INVX4 U708 ( .IN(n844), .OUT(n865) );
  NOR2X1 U709 ( .IN1(n1058), .IN2(StateMC[1]), .OUT(n827) );
  NOR2X1 U710 ( .IN1(n851), .IN2(Adder_ack), .OUT(n286) );
  NANDX2 U711 ( .IN1(n285), .IN2(n825), .OUT(n1130) );
  NOR2X1 U712 ( .IN1(RSTn_BAR), .IN2(n1138), .OUT(n569) );
  AOI22 U713 ( .IN1(n288), .IN2(n230), .IN3(Adder_dataout[8]), .IN4(n569), 
        .OUT(n289) );
  NOR2X1 U714 ( .IN1(n290), .IN2(StateMC[1]), .OUT(n824) );
  NANDX2 U715 ( .IN1(n285), .IN2(n824), .OUT(n1146) );
  OAI21 U716 ( .IN1(StateMC[0]), .IN2(n870), .IN3(n285), .OUT(n579) );
  NANDX2 U717 ( .IN1(n885), .IN2(n886), .OUT(n1116) );
  AOI22 U718 ( .IN1(Op2_Sign_reg), .IN2(n1052), .IN3(Datain1[15]), .IN4(n821), 
        .OUT(n292) );
  OAI21 U719 ( .IN1(n1116), .IN2(n293), .IN3(n292), .OUT(n1090) );
  AOI22 U720 ( .IN1(Op1_Sign_reg), .IN2(n1052), .IN3(Datain2[15]), .IN4(n821), 
        .OUT(n294) );
  OAI21 U721 ( .IN1(n1116), .IN2(n295), .IN3(n294), .OUT(n1081) );
  INVX4 U722 ( .IN(n815), .OUT(n727) );
  NOR2X1 U723 ( .IN1(n276), .IN2(n304), .OUT(n301) );
  NOR2X1 U724 ( .IN1(n281), .IN2(n280), .OUT(n300) );
  NOR2X1 U725 ( .IN1(n279), .IN2(n237), .OUT(n303) );
  NOR2X1 U726 ( .IN1(n233), .IN2(n304), .OUT(n305) );
  NAND3X1 U727 ( .IN1(n757), .IN2(n608), .IN3(n601), .OUT(n307) );
  NOR2X1 U728 ( .IN1(n275), .IN2(n208), .OUT(n309) );
  NOR2X1 U729 ( .IN1(n284), .IN2(n275), .OUT(n311) );
  NAND3X1 U730 ( .IN1(n764), .IN2(n594), .IN3(n669), .OUT(n804) );
  NOR2X1 U731 ( .IN1(n739), .IN2(n804), .OUT(n315) );
  AOI22 U732 ( .IN1(n474), .IN2(n283), .IN3(n275), .IN4(n450), .OUT(n324) );
  AOI22 U733 ( .IN1(n473), .IN2(n284), .IN3(n276), .IN4(n546), .OUT(n323) );
  NOR2X1 U734 ( .IN1(n283), .IN2(n282), .OUT(n334) );
  MUX2X1 U735 ( .IN1(n233), .IN2(n276), .S(n345), .OUT(n359) );
  AOI22 U736 ( .IN1(n210), .IN2(n276), .IN3(n275), .IN4(n233), .OUT(n330) );
  AOI22 U737 ( .IN1(n826), .IN2(Adder_dataout[1]), .IN3(n278), .IN4(n537), 
        .OUT(n329) );
  OAI21 U738 ( .IN1(n330), .IN2(n535), .IN3(n329), .OUT(n331) );
  AOI21 U739 ( .IN1(n526), .IN2(n445), .IN3(n331), .OUT(n332) );
  OAI21 U740 ( .IN1(n516), .IN2(n333), .IN3(n332), .OUT(n379) );
  OAI21 U741 ( .IN1(n284), .IN2(n358), .IN3(n275), .OUT(n335) );
  NOR2X1 U742 ( .IN1(n281), .IN2(Final_Mantissa_reg[9]), .OUT(n337) );
  NOR2X1 U743 ( .IN1(n282), .IN2(n278), .OUT(n336) );
  MUX2X1 U744 ( .IN1(n280), .IN2(n231), .S(n339), .OUT(n480) );
  MUX2X1 U745 ( .IN1(n281), .IN2(n209), .S(n340), .OUT(n485) );
  NOR2X1 U746 ( .IN1(n480), .IN2(n485), .OUT(n343) );
  MUX2X1 U747 ( .IN1(n232), .IN2(Final_Mantissa_reg[9]), .S(n342), .OUT(n471)
         );
  NOR2X1 U748 ( .IN1(n387), .IN2(n748), .OUT(n352) );
  MUX2X1 U749 ( .IN1(n279), .IN2(n206), .S(n347), .OUT(n481) );
  OAI21 U750 ( .IN1(n276), .IN2(n345), .IN3(n278), .OUT(n346) );
  NOR2X1 U751 ( .IN1(n481), .IN2(n398), .OUT(n349) );
  NAND3X1 U752 ( .IN1(n350), .IN2(n398), .IN3(n445), .OUT(n351) );
  NOR2X1 U753 ( .IN1(n354), .IN2(n556), .OUT(n355) );
  NAND3X1 U754 ( .IN1(n636), .IN2(n755), .IN3(n621), .OUT(n363) );
  MUX2X1 U755 ( .IN1(n208), .IN2(n284), .S(n358), .OUT(n382) );
  NAND3X1 U756 ( .IN1(n387), .IN2(n398), .IN3(n359), .OUT(n361) );
  NOR2X1 U757 ( .IN1(n363), .IN2(n656), .OUT(n364) );
  NAND3X1 U758 ( .IN1(n662), .IN2(n266), .IN3(n621), .OUT(n368) );
  NAND3X1 U759 ( .IN1(n282), .IN2(n283), .IN3(n284), .OUT(n365) );
  NOR2X1 U760 ( .IN1(n368), .IN2(n654), .OUT(n369) );
  INVX4 U761 ( .IN(n505), .OUT(n484) );
  INVX4 U762 ( .IN(n722), .OUT(n750) );
  NOR2X1 U763 ( .IN1(n382), .IN2(n373), .OUT(n772) );
  NOR2X1 U764 ( .IN1(n374), .IN2(n772), .OUT(n400) );
  AOI22 U765 ( .IN1(n546), .IN2(n477), .IN3(n484), .IN4(n439), .OUT(n377) );
  NOR2X1 U766 ( .IN1(n236), .IN2(n377), .OUT(n378) );
  OAI21 U767 ( .IN1(n379), .IN2(n378), .IN3(n285), .OUT(n391) );
  NOR2X1 U768 ( .IN1(StateMC[0]), .IN2(n897), .OUT(n1145) );
  NOR2X1 U769 ( .IN1(n825), .IN2(n1145), .OUT(n820) );
  AOI21 U770 ( .IN1(n220), .IN2(StateMC[2]), .IN3(RSTn_BAR), .OUT(n715) );
  OAI21 U771 ( .IN1(RSTn_BAR), .IN2(n539), .IN3(n567), .OUT(n518) );
  AOI22 U772 ( .IN1(n482), .IN2(n490), .IN3(n525), .IN4(n479), .OUT(n389) );
  AOI22 U773 ( .IN1(n486), .IN2(n513), .IN3(n484), .IN4(n445), .OUT(n388) );
  AOI22 U774 ( .IN1(n276), .IN2(n518), .IN3(n417), .IN4(n487), .OUT(n390) );
  AOI22 U775 ( .IN1(n479), .IN2(n282), .IN3(n484), .IN4(n525), .OUT(n392) );
  AOI22 U776 ( .IN1(n450), .IN2(n283), .IN3(n546), .IN4(n284), .OUT(n396) );
  NOR2X1 U777 ( .IN1(n722), .IN2(n400), .OUT(n803) );
  NOR2X1 U778 ( .IN1(n847), .IN2(n505), .OUT(n401) );
  AOI22 U779 ( .IN1(n546), .IN2(n472), .IN3(n803), .IN4(n401), .OUT(n415) );
  NAND3X1 U780 ( .IN1(n539), .IN2(n405), .IN3(n502), .OUT(n478) );
  AOI22 U781 ( .IN1(n826), .IN2(Adder_dataout[5]), .IN3(Final_Mantissa_reg[9]), 
        .IN4(n537), .OUT(n404) );
  OAI21 U782 ( .IN1(n405), .IN2(n430), .IN3(n404), .OUT(n406) );
  AOI21 U783 ( .IN1(n526), .IN2(n485), .IN3(n406), .OUT(n412) );
  AOI22 U784 ( .IN1(n474), .IN2(n278), .IN3(n279), .IN4(n473), .OUT(n407) );
  OAI21 U785 ( .IN1(n231), .IN2(n475), .IN3(n407), .OUT(n408) );
  NAND3X1 U786 ( .IN1(n412), .IN2(n411), .IN3(n410), .OUT(n413) );
  AOI21 U787 ( .IN1(n478), .IN2(n281), .IN3(n413), .OUT(n414) );
  OAI21 U788 ( .IN1(n236), .IN2(n415), .IN3(n414), .OUT(n416) );
  AOI21 U789 ( .IN1(n439), .IN2(n417), .IN3(n416), .OUT(n422) );
  AOI22 U790 ( .IN1(n456), .IN2(n482), .IN3(n481), .IN4(n479), .OUT(n419) );
  AOI22 U791 ( .IN1(n486), .IN2(n480), .IN3(n484), .IN4(n485), .OUT(n418) );
  AOI22 U792 ( .IN1(n281), .IN2(n561), .IN3(n420), .IN4(n487), .OUT(n421) );
  OAI21 U793 ( .IN1(RSTn_BAR), .IN2(n422), .IN3(n421), .OUT(n1064) );
  AOI22 U794 ( .IN1(n482), .IN2(n282), .IN3(n490), .IN4(n479), .OUT(n424) );
  AOI22 U795 ( .IN1(n486), .IN2(n525), .IN3(n513), .IN4(n484), .OUT(n423) );
  AOI22 U796 ( .IN1(n282), .IN2(n474), .IN3(n284), .IN4(n450), .OUT(n426) );
  AOI22 U797 ( .IN1(n473), .IN2(n283), .IN3(n275), .IN4(n546), .OUT(n425) );
  AOI22 U798 ( .IN1(n474), .IN2(n276), .IN3(n279), .IN4(n450), .OUT(n428) );
  AOI22 U799 ( .IN1(n473), .IN2(n278), .IN3(n280), .IN4(n546), .OUT(n427) );
  AOI21 U800 ( .IN1(n510), .IN2(n739), .IN3(n429), .OUT(n436) );
  OAI21 U801 ( .IN1(n280), .IN2(n431), .IN3(n430), .OUT(n433) );
  AOI22 U802 ( .IN1(n826), .IN2(Adder_dataout[4]), .IN3(n281), .IN4(n537), 
        .OUT(n432) );
  OAI21 U803 ( .IN1(n535), .IN2(n433), .IN3(n432), .OUT(n434) );
  AOI21 U804 ( .IN1(n526), .IN2(n480), .IN3(n434), .OUT(n435) );
  OAI21 U805 ( .IN1(n437), .IN2(n436), .IN3(n435), .OUT(n438) );
  AOI21 U806 ( .IN1(n439), .IN2(n509), .IN3(n438), .OUT(n444) );
  AOI22 U807 ( .IN1(n482), .IN2(n445), .IN3(n456), .IN4(n479), .OUT(n441) );
  AOI22 U808 ( .IN1(n486), .IN2(n481), .IN3(n484), .IN4(n480), .OUT(n440) );
  AOI22 U809 ( .IN1(n280), .IN2(n518), .IN3(n442), .IN4(n487), .OUT(n443) );
  OAI21 U810 ( .IN1(RSTn_BAR), .IN2(n444), .IN3(n443), .OUT(n1065) );
  AOI22 U811 ( .IN1(n482), .IN2(n525), .IN3(n513), .IN4(n479), .OUT(n447) );
  AOI22 U812 ( .IN1(n486), .IN2(n445), .IN3(n456), .IN4(n484), .OUT(n446) );
  AOI22 U813 ( .IN1(n486), .IN2(n282), .IN3(n484), .IN4(n490), .OUT(n465) );
  AOI22 U814 ( .IN1(n284), .IN2(n474), .IN3(n276), .IN4(n450), .OUT(n449) );
  AOI22 U815 ( .IN1(n473), .IN2(n275), .IN3(n278), .IN4(n546), .OUT(n448) );
  AOI22 U816 ( .IN1(n450), .IN2(n282), .IN3(n283), .IN4(n546), .OUT(n458) );
  OAI21 U817 ( .IN1(n278), .IN2(n452), .IN3(n451), .OUT(n454) );
  AOI22 U818 ( .IN1(n826), .IN2(Adder_dataout[2]), .IN3(n279), .IN4(n537), 
        .OUT(n453) );
  OAI21 U819 ( .IN1(n535), .IN2(n454), .IN3(n453), .OUT(n455) );
  AOI21 U820 ( .IN1(n456), .IN2(n526), .IN3(n455), .OUT(n457) );
  OAI21 U821 ( .IN1(n459), .IN2(n458), .IN3(n457), .OUT(n460) );
  AOI21 U822 ( .IN1(n527), .IN2(n476), .IN3(n460), .OUT(n461) );
  OAI21 U823 ( .IN1(n465), .IN2(n558), .IN3(n461), .OUT(n462) );
  AOI21 U824 ( .IN1(n554), .IN2(n467), .IN3(n462), .OUT(n464) );
  OAI21 U825 ( .IN1(RSTn_BAR), .IN2(n464), .IN3(n463), .OUT(n1067) );
  NOR2X1 U826 ( .IN1(n466), .IN2(n465), .OUT(n493) );
  MUX2X1 U827 ( .IN1(n283), .IN2(n282), .S(n718), .OUT(n469) );
  NOR2X1 U828 ( .IN1(n739), .IN2(n769), .OUT(n468) );
  AOI22 U829 ( .IN1(n826), .IN2(n240), .IN3(n283), .IN4(n565), .OUT(n488) );
  OAI21 U830 ( .IN1(n208), .IN2(n523), .IN3(n488), .OUT(n489) );
  AOI21 U831 ( .IN1(n526), .IN2(n490), .IN3(n489), .OUT(n497) );
  NAND3X1 U832 ( .IN1(n492), .IN2(n745), .IN3(n491), .OUT(n496) );
  NAND3X1 U833 ( .IN1(n497), .IN2(n496), .IN3(n495), .OUT(n498) );
  AOI22 U834 ( .IN1(n283), .IN2(n533), .IN3(n285), .IN4(n498), .OUT(n672) );
  NAND3X1 U835 ( .IN1(n1105), .IN2(n1104), .IN3(n1146), .OUT(n732) );
  OAI21 U836 ( .IN1(n732), .IN2(n817), .IN3(n211), .OUT(n500) );
  NOR2X1 U837 ( .IN1(RSTn_BAR), .IN2(n238), .OUT(n501) );
  AOI22 U838 ( .IN1(n569), .IN2(n211), .IN3(n501), .IN4(n537), .OUT(n508) );
  NAND3X1 U839 ( .IN1(n820), .IN2(n545), .IN3(n502), .OUT(n503) );
  AOI21 U840 ( .IN1(n503), .IN2(n285), .IN3(n533), .OUT(n504) );
  OAI21 U841 ( .IN1(n505), .IN2(n520), .IN3(n504), .OUT(n506) );
  AOI22 U842 ( .IN1(n826), .IN2(Adder_dataout[0]), .IN3(n276), .IN4(n537), 
        .OUT(n511) );
  OAI21 U843 ( .IN1(n275), .IN2(n535), .IN3(n511), .OUT(n512) );
  AOI21 U844 ( .IN1(n526), .IN2(n513), .IN3(n512), .OUT(n514) );
  OAI21 U845 ( .IN1(n516), .IN2(n515), .IN3(n514), .OUT(n517) );
  AOI22 U846 ( .IN1(n275), .IN2(n518), .IN3(n285), .IN4(n517), .OUT(n519) );
  OAI21 U847 ( .IN1(n521), .IN2(n520), .IN3(n519), .OUT(n1069) );
  AOI22 U848 ( .IN1(n826), .IN2(n226), .IN3(n284), .IN4(n565), .OUT(n522) );
  OAI21 U849 ( .IN1(n210), .IN2(n523), .IN3(n522), .OUT(n524) );
  AOI21 U850 ( .IN1(n526), .IN2(n525), .IN3(n524), .OUT(n531) );
  NAND3X1 U851 ( .IN1(n531), .IN2(n530), .IN3(n529), .OUT(n532) );
  AOI22 U852 ( .IN1(n284), .IN2(n533), .IN3(n285), .IN4(n532), .OUT(n664) );
  NOR2X1 U853 ( .IN1(n534), .IN2(n536), .OUT(n563) );
  NOR2X1 U854 ( .IN1(n535), .IN2(n563), .OUT(n542) );
  OAI21 U855 ( .IN1(n232), .IN2(n536), .IN3(n205), .OUT(n541) );
  AOI22 U856 ( .IN1(n826), .IN2(Adder_dataout[7]), .IN3(carry_reg), .IN4(n537), 
        .OUT(n538) );
  OAI21 U857 ( .IN1(n205), .IN2(n539), .IN3(n538), .OUT(n540) );
  AOI21 U858 ( .IN1(n542), .IN2(n541), .IN3(n540), .OUT(n543) );
  OAI21 U859 ( .IN1(n545), .IN2(n544), .IN3(n543), .OUT(n553) );
  NOR2X1 U860 ( .IN1(Final_Mantissa_reg[10]), .IN2(n739), .OUT(n547) );
  OAI21 U861 ( .IN1(n549), .IN2(n548), .IN3(n805), .OUT(n550) );
  AOI21 U862 ( .IN1(n551), .IN2(n550), .IN3(n847), .OUT(n552) );
  NOR2X1 U863 ( .IN1(n553), .IN2(n552), .OUT(n559) );
  OAI21 U864 ( .IN1(n556), .IN2(n555), .IN3(n554), .OUT(n557) );
  NAND3X1 U865 ( .IN1(n559), .IN2(n558), .IN3(n557), .OUT(n560) );
  AOI22 U866 ( .IN1(n561), .IN2(Final_Mantissa_reg[10]), .IN3(n285), .IN4(n560), .OUT(n562) );
  NAND3X1 U867 ( .IN1(n1146), .IN2(n567), .IN3(n566), .OUT(n568) );
  AOI22 U868 ( .IN1(n569), .IN2(Adder_carryout), .IN3(carry_reg), .IN4(n568), 
        .OUT(n570) );
  OAI21 U869 ( .IN1(n717), .IN2(n1125), .IN3(n570), .OUT(n1061) );
  INVX4 U870 ( .IN(n1146), .OUT(n823) );
  NOR2X1 U871 ( .IN1(n572), .IN2(n571), .OUT(n576) );
  NOR2X1 U872 ( .IN1(n574), .IN2(n573), .OUT(n575) );
  OAI21 U873 ( .IN1(n750), .IN2(n696), .IN3(n823), .OUT(n583) );
  INVX4 U874 ( .IN(n583), .OUT(n650) );
  AOI22 U875 ( .IN1(DP_OP_986_157_3518_n93), .IN2(n647), .IN3(Datain1[10]), 
        .IN4(n822), .OUT(n586) );
  NAND3X1 U876 ( .IN1(n586), .IN2(n585), .IN3(n584), .OUT(n1097) );
  NOR2X1 U877 ( .IN1(Final_Exponent_reg[6]), .IN2(n145), .OUT(n588) );
  NOR2X1 U878 ( .IN1(Final_Exponent_reg[4]), .IN2(Final_Exponent_reg[7]), 
        .OUT(n587) );
  AOI22 U879 ( .IN1(n692), .IN2(n805), .IN3(n750), .IN4(n772), .OUT(n597) );
  OAI21 U880 ( .IN1(Final_Exponent_reg[1]), .IN2(Final_Exponent_reg[2]), .IN3(
        DP_OP_986_157_3518_n93), .OUT(n592) );
  OAI21 U881 ( .IN1(n722), .IN2(n754), .IN3(n595), .OUT(n596) );
  OAI21 U882 ( .IN1(n691), .IN2(n597), .IN3(n644), .OUT(n599) );
  AOI22 U883 ( .IN1(n598), .IN2(n805), .IN3(n750), .IN4(n654), .OUT(n703) );
  NOR2X1 U884 ( .IN1(n653), .IN2(n703), .OUT(n627) );
  NOR2X1 U885 ( .IN1(n599), .IN2(n627), .OUT(n600) );
  AOI22 U886 ( .IN1(n759), .IN2(n805), .IN3(n750), .IN4(n752), .OUT(n605) );
  OAI21 U887 ( .IN1(Final_Exponent_reg[0]), .IN2(n606), .IN3(n607), .OUT(n684)
         );
  NOR2X1 U888 ( .IN1(n757), .IN2(n684), .OUT(n604) );
  NOR2X1 U889 ( .IN1(n722), .IN2(n684), .OUT(n603) );
  AOI22 U890 ( .IN1(n604), .IN2(n805), .IN3(n603), .IN4(n665), .OUT(n637) );
  OAI21 U891 ( .IN1(n674), .IN2(n605), .IN3(n637), .OUT(n615) );
  AOI22 U892 ( .IN1(n673), .IN2(n805), .IN3(n750), .IN4(n659), .OUT(n609) );
  OAI21 U893 ( .IN1(n722), .IN2(n657), .IN3(n613), .OUT(n614) );
  NOR2X1 U894 ( .IN1(n615), .IN2(n617), .OUT(n616) );
  NAND3X1 U895 ( .IN1(n682), .IN2(n663), .IN3(n805), .OUT(n626) );
  NAND3X1 U896 ( .IN1(n750), .IN2(n663), .IN3(n619), .OUT(n625) );
  NOR2X1 U897 ( .IN1(n675), .IN2(n646), .OUT(n623) );
  NOR2X1 U898 ( .IN1(n722), .IN2(n676), .OUT(n622) );
  AOI22 U899 ( .IN1(n624), .IN2(n623), .IN3(n622), .IN4(n658), .OUT(n640) );
  NAND3X1 U900 ( .IN1(n626), .IN2(n625), .IN3(n640), .OUT(n628) );
  NOR2X1 U901 ( .IN1(n628), .IN2(n627), .OUT(n629) );
  OAI21 U902 ( .IN1(n762), .IN2(n632), .IN3(n707), .OUT(n633) );
  AOI21 U903 ( .IN1(n635), .IN2(n634), .IN3(n633), .OUT(n639) );
  NAND3X1 U904 ( .IN1(n750), .IN2(n660), .IN3(n661), .OUT(n638) );
  NAND3X1 U905 ( .IN1(n639), .IN2(n638), .IN3(n637), .OUT(n642) );
  NOR2X1 U906 ( .IN1(n642), .IN2(n641), .OUT(n645) );
  NAND3X1 U907 ( .IN1(n645), .IN2(n644), .IN3(n643), .OUT(C1_Z_0) );
  AOI22 U908 ( .IN1(Final_Exponent_reg[7]), .IN2(n647), .IN3(Datain1[14]), 
        .IN4(n822), .OUT(n648) );
  AOI21 U909 ( .IN1(n821), .IN2(DP_OP_982J1_125_6202_n102), .IN3(n649), .OUT(
        n652) );
  AOI21 U910 ( .IN1(n654), .IN2(n653), .IN3(n722), .OUT(n668) );
  OAI21 U911 ( .IN1(n704), .IN2(n669), .IN3(n805), .OUT(n670) );
  AOI22 U912 ( .IN1(n674), .IN2(n759), .IN3(n673), .IN4(n671), .OUT(n679) );
  AOI22 U913 ( .IN1(n684), .IN2(n683), .IN3(n682), .IN4(n681), .OUT(n688) );
  NAND3X1 U914 ( .IN1(n689), .IN2(n688), .IN3(n687), .OUT(n698) );
  AOI22 U915 ( .IN1(n692), .IN2(n691), .IN3(n690), .IN4(n761), .OUT(n693) );
  OAI21 U916 ( .IN1(n695), .IN2(n694), .IN3(n693), .OUT(n699) );
  NAND3X1 U917 ( .IN1(n722), .IN2(n740), .IN3(n697), .OUT(n701) );
  NOR2X1 U918 ( .IN1(n699), .IN2(n698), .OUT(n711) );
  AOI22 U919 ( .IN1(exc_reg_0_), .IN2(n701), .IN3(n805), .IN4(n700), .OUT(n702) );
  OAI21 U920 ( .IN1(n704), .IN2(n703), .IN3(n702), .OUT(n705) );
  AOI21 U921 ( .IN1(n706), .IN2(n750), .IN3(n705), .OUT(n714) );
  AOI21 U922 ( .IN1(n711), .IN2(n710), .IN3(n709), .OUT(n712) );
  AOI21 U923 ( .IN1(n836), .IN2(n712), .IN3(n222), .OUT(n725) );
  MUX2X1 U924 ( .IN1(n725), .IN2(n819), .S(n714), .OUT(n838) );
  AOI22 U925 ( .IN1(Final_Mantissa_reg[10]), .IN2(n719), .IN3(n805), .IN4(n718), .OUT(n720) );
  OAI21 U926 ( .IN1(n722), .IN2(n721), .IN3(n720), .OUT(n723) );
  AOI22 U927 ( .IN1(Debug_reg[0]), .IN2(n1144), .IN3(n823), .IN4(n723), .OUT(
        n724) );
  AOI22 U928 ( .IN1(Exc_value[2]), .IN2(n893), .IN3(n823), .IN4(n725), .OUT(
        n890) );
  NAND3X1 U929 ( .IN1(n727), .IN2(n204), .IN3(n726), .OUT(n728) );
  NAND3X1 U930 ( .IN1(n1058), .IN2(n1138), .IN3(n728), .OUT(n1059) );
  AOI22 U931 ( .IN1(n732), .IN2(n226), .IN3(n1106), .IN4(n817), .OUT(n1107) );
  AOI21 U932 ( .IN1(n211), .IN2(n240), .IN3(n729), .OUT(n731) );
  OAI21 U933 ( .IN1(add_x_35_A_0_), .IN2(n729), .IN3(add_x_35_A_1_), .OUT(n730) );
  OAI21 U934 ( .IN1(n732), .IN2(n731), .IN3(n730), .OUT(n1123) );
  AOI21 U935 ( .IN1(n734), .IN2(Op1_Sign_reg), .IN3(n733), .OUT(n1127) );
  NOR2X1 U936 ( .IN1(n277), .IN2(RSTn_BAR), .OUT(n735) );
  AOI22 U937 ( .IN1(n1144), .IN2(n251), .IN3(n737), .IN4(n750), .OUT(n1126) );
  NOR2X1 U938 ( .IN1(n738), .IN2(n762), .OUT(n744) );
  OAI21 U939 ( .IN1(n742), .IN2(n741), .IN3(n740), .OUT(n743) );
  AOI21 U940 ( .IN1(n745), .IN2(n744), .IN3(n743), .OUT(n746) );
  OAI21 U941 ( .IN1(n748), .IN2(n747), .IN3(n746), .OUT(n1140) );
  NAND3X1 U942 ( .IN1(n751), .IN2(n750), .IN3(n749), .OUT(n753) );
  NOR2X1 U943 ( .IN1(n753), .IN2(n752), .OUT(n756) );
  NAND3X1 U944 ( .IN1(n756), .IN2(n755), .IN3(n754), .OUT(n771) );
  NAND3X1 U945 ( .IN1(n758), .IN2(n277), .IN3(n757), .OUT(n760) );
  NOR2X1 U946 ( .IN1(n760), .IN2(n759), .OUT(n765) );
  NOR2X1 U947 ( .IN1(n762), .IN2(n761), .OUT(n763) );
  NAND3X1 U948 ( .IN1(n765), .IN2(n764), .IN3(n763), .OUT(n766) );
  AOI21 U949 ( .IN1(n805), .IN2(n769), .IN3(n768), .OUT(n770) );
  OAI21 U950 ( .IN1(n772), .IN2(n771), .IN3(n770), .OUT(n1142) );
  AOI22 U951 ( .IN1(n272), .IN2(n250), .IN3(n275), .IN4(n865), .OUT(n773) );
  AOI22 U952 ( .IN1(n272), .IN2(n225), .IN3(n276), .IN4(n865), .OUT(n774) );
  AOI22 U953 ( .IN1(n272), .IN2(n249), .IN3(n278), .IN4(n865), .OUT(n775) );
  AOI22 U954 ( .IN1(n272), .IN2(n221), .IN3(n279), .IN4(n865), .OUT(n776) );
  AOI22 U955 ( .IN1(n272), .IN2(n248), .IN3(n280), .IN4(n865), .OUT(n777) );
  AOI22 U956 ( .IN1(n272), .IN2(n224), .IN3(n281), .IN4(n865), .OUT(n778) );
  AOI22 U957 ( .IN1(n272), .IN2(n247), .IN3(Final_Mantissa_reg[9]), .IN4(n865), 
        .OUT(n779) );
  AOI22 U958 ( .IN1(n272), .IN2(Op2_Mantissa_reg_7_), .IN3(
        Final_Exponent_reg[0]), .IN4(n865), .OUT(ExcCheck_Datain_7__BAR) );
  AOI22 U959 ( .IN1(Final_Exponent_reg[0]), .IN2(n272), .IN3(
        Final_Exponent_reg[1]), .IN4(n865), .OUT(n781) );
  AOI22 U960 ( .IN1(Final_Exponent_reg[1]), .IN2(n272), .IN3(
        Final_Exponent_reg[2]), .IN4(n865), .OUT(n782) );
  AOI22 U961 ( .IN1(Final_Exponent_reg[2]), .IN2(n272), .IN3(
        DP_OP_986_157_3518_n93), .IN4(n865), .OUT(ExcCheck_Datain_10__BAR) );
  AOI22 U962 ( .IN1(DP_OP_986_157_3518_n93), .IN2(n272), .IN3(
        Final_Exponent_reg[4]), .IN4(n865), .OUT(n784) );
  AOI22 U963 ( .IN1(Final_Exponent_reg[4]), .IN2(n272), .IN3(n145), .IN4(n865), 
        .OUT(n785) );
  AOI22 U964 ( .IN1(n145), .IN2(n272), .IN3(Final_Exponent_reg[6]), .IN4(n865), 
        .OUT(ExcCheck_Datain_13__BAR) );
  AOI22 U965 ( .IN1(Final_Exponent_reg[6]), .IN2(n272), .IN3(
        Final_Exponent_reg[7]), .IN4(n865), .OUT(n786) );
  INVX4 U966 ( .IN(n862), .OUT(n800) );
  AOI21 U967 ( .IN1(n805), .IN2(n804), .IN3(n803), .OUT(n806) );
  OAI21 U968 ( .IN1(n1146), .IN2(n806), .IN3(n1139), .OUT(n112) );
  MUX2X1 U969 ( .IN1(n247), .IN2(add_x_35_A_9_), .S(n807), .OUT(n808) );
  NOR2X1 U970 ( .IN1(n1130), .IN2(n808), .OUT(n122) );
  MUX2X1 U971 ( .IN1(n248), .IN2(add_x_35_A_7_), .S(n809), .OUT(n810) );
  NOR2X1 U972 ( .IN1(n1130), .IN2(n810), .OUT(n120) );
  MUX2X1 U973 ( .IN1(n249), .IN2(add_x_35_A_5_), .S(n811), .OUT(n812) );
  NOR2X1 U974 ( .IN1(n1130), .IN2(n812), .OUT(n118) );
  MUX2X1 U975 ( .IN1(n250), .IN2(add_x_35_A_3_), .S(n813), .OUT(n814) );
  NOR2X1 U976 ( .IN1(n1130), .IN2(n814), .OUT(n116) );
  OAI21 U977 ( .IN1(Op2_Mantissa_reg_7_), .IN2(n816), .IN3(n817), .OUT(n818)
         );
  NOR2X1 U978 ( .IN1(StateMC[0]), .IN2(n204), .OUT(n840) );
  NOR2X1 U979 ( .IN1(n241), .IN2(n846), .OUT(n866) );
  INVX1 U980 ( .IN(Exc_value[1]), .OUT(n830) );
  INVX1 U981 ( .IN(Exc_value[2]), .OUT(n828) );
  AOI22 U982 ( .IN1(Exc_value[2]), .IN2(Exc_value[0]), .IN3(n830), .IN4(n828), 
        .OUT(n829) );
  AOI21 U983 ( .IN1(Exc_value[0]), .IN2(n830), .IN3(n829), .OUT(n832) );
  NOR2X1 U984 ( .IN1(n827), .IN2(n826), .OUT(n831) );
  OAI21 U985 ( .IN1(n835), .IN2(n832), .IN3(n831), .OUT(n833) );
  OAI21 U986 ( .IN1(n840), .IN2(n833), .IN3(n285), .OUT(n915) );
  AOI22 U987 ( .IN1(n223), .IN2(n222), .IN3(exc_reg_0_), .IN4(n242), .OUT(n834) );
  AOI21 U988 ( .IN1(n222), .IN2(exc_reg_0_), .IN3(n834), .OUT(n861) );
  OAI21 U989 ( .IN1(n861), .IN2(n1138), .IN3(n835), .OUT(n850) );
  NAND2X1 U990 ( .IN1(n838), .IN2(n837), .OUT(n839) );
  AOI22 U991 ( .IN1(n827), .IN2(n1125), .IN3(n824), .IN4(n839), .OUT(n841) );
  NAND2X1 U992 ( .IN1(StateMC[1]), .IN2(n840), .OUT(n844) );
  NAND3X1 U993 ( .IN1(n820), .IN2(n841), .IN3(n844), .OUT(n842) );
  OAI21 U994 ( .IN1(n850), .IN2(n842), .IN3(n285), .OUT(n922) );
  NOR2X1 U995 ( .IN1(n272), .IN2(n825), .OUT(n843) );
  AOI22 U996 ( .IN1(StateMC[0]), .IN2(n845), .IN3(n865), .IN4(Exc_Ack), .OUT(
        n848) );
  NOR2X1 U997 ( .IN1(StateMC[0]), .IN2(n846), .OUT(n868) );
  NAND3X1 U998 ( .IN1(n848), .IN2(n884), .IN3(n847), .OUT(n849) );
  OAI21 U999 ( .IN1(n850), .IN2(n849), .IN3(n285), .OUT(n991) );
  NOR2X1 U1000 ( .IN1(n204), .IN2(n851), .OUT(Dataout_valid) );
  NOR2X1 U1001 ( .IN1(n274), .IN2(n862), .OUT(Dataout[15]) );
  INVX1 U1002 ( .IN(Mode[1]), .OUT(n853) );
  NAND2X1 U1003 ( .IN1(Mode[0]), .IN2(n853), .OUT(n852) );
  NOR2X1 U1004 ( .IN1(Mode[2]), .IN2(n852), .OUT(n858) );
  NOR2X1 U1005 ( .IN1(Mode[2]), .IN2(n853), .OUT(n859) );
  AOI22 U1006 ( .IN1(StateMC[0]), .IN2(n858), .IN3(Debug_reg[0]), .IN4(n859), 
        .OUT(n854) );
  AOI22 U1007 ( .IN1(StateMC[1]), .IN2(n858), .IN3(Debug_reg[1]), .IN4(n859), 
        .OUT(n855) );
  AOI22 U1008 ( .IN1(StateMC[2]), .IN2(n858), .IN3(Debug_reg[2]), .IN4(n859), 
        .OUT(n856) );
  NAND2X1 U1009 ( .IN1(Debug_reg[3]), .IN2(n859), .OUT(n857) );
  AOI21 U1010 ( .IN1(n859), .IN2(Debug_valid_reg), .IN3(n858), .OUT(n860) );
  NOR2X1 U1011 ( .IN1(n862), .IN2(n861), .OUT(n863) );
  NOR2X1 U1012 ( .IN1(n243), .IN2(n864), .OUT(Exc[0]) );
  NOR2X1 U1013 ( .IN1(n223), .IN2(n864), .OUT(Exc[1]) );
  NOR2X1 U1014 ( .IN1(n222), .IN2(n864), .OUT(Exc[2]) );
  NOR2X1 U1015 ( .IN1(n219), .IN2(n1130), .OUT(N252) );
  NOR2X1 U1016 ( .IN1(n218), .IN2(n1130), .OUT(N253) );
  NOR2X1 U1017 ( .IN1(n217), .IN2(n1130), .OUT(N254) );
  NOR2X1 U1018 ( .IN1(n216), .IN2(n1130), .OUT(N255) );
  NOR2X1 U1019 ( .IN1(n215), .IN2(n1130), .OUT(N256) );
  NOR2X1 U1020 ( .IN1(n214), .IN2(n1130), .OUT(N257) );
  NOR2X1 U1021 ( .IN1(n213), .IN2(n1130), .OUT(N258) );
  NOR2X1 U1022 ( .IN1(n212), .IN2(n1130), .OUT(N259) );
  OAI21 U1023 ( .IN1(n272), .IN2(n865), .IN3(n285), .OUT(n1104) );
  NOR2X1 U1024 ( .IN1(Exc_Ack), .IN2(n1104), .OUT(N270) );
  INVX1 U1025 ( .IN(Data_valid), .OUT(n867) );
  AOI21 U1026 ( .IN1(DP_OP_982J1_125_6202_n102), .IN2(n906), .IN3(
        DP_OP_982J1_125_6202_n101), .OUT(n882) );
  AOI22 U1027 ( .IN1(DP_OP_982J1_125_6202_n100), .IN2(n199), .IN3(
        DP_OP_982J1_125_6202_n101), .IN4(n200), .OUT(n881) );
  AOI22 U1028 ( .IN1(DP_OP_982J1_125_6202_n91), .IN2(n179), .IN3(Datain1[12]), 
        .IN4(n144), .OUT(n879) );
  AOI22 U1029 ( .IN1(Datain2[7]), .IN2(n181), .IN3(Datain2[8]), .IN4(n194), 
        .OUT(n871) );
  AOI21 U1030 ( .IN1(Datain1[8]), .IN2(n176), .IN3(n871), .OUT(n873) );
  NOR2X1 U1031 ( .IN1(n873), .IN2(DP_OP_982J1_125_6202_n97), .OUT(n875) );
  NOR2X1 U1032 ( .IN1(Datain1[10]), .IN2(n178), .OUT(n872) );
  AOI21 U1033 ( .IN1(DP_OP_982J1_125_6202_n97), .IN2(n873), .IN3(n872), .OUT(
        n874) );
  OAI21 U1034 ( .IN1(Datain1[9]), .IN2(n875), .IN3(n874), .OUT(n876) );
  OAI21 U1035 ( .IN1(Datain2[10]), .IN2(n196), .IN3(n876), .OUT(n877) );
  OAI21 U1036 ( .IN1(DP_OP_982J1_125_6202_n91), .IN2(n179), .IN3(n877), .OUT(
        n878) );
  AOI22 U1037 ( .IN1(DP_OP_982J1_125_6202_n102), .IN2(n906), .IN3(n879), .IN4(
        n878), .OUT(n880) );
  AOI22 U1038 ( .IN1(Datain1[13]), .IN2(n882), .IN3(n881), .IN4(n880), .OUT(
        n883) );
  OAI21 U1039 ( .IN1(DP_OP_982J1_125_6202_n102), .IN2(n906), .IN3(n883), .OUT(
        n886) );
  NOR2X1 U1040 ( .IN1(n884), .IN2(RSTn_BAR), .OUT(n885) );
  MUX2X1 U1041 ( .IN1(n220), .IN2(n241), .S(StateMC[2]), .OUT(n887) );
  NOR2X1 U1042 ( .IN1(n887), .IN2(RSTn_BAR), .OUT(n888) );
  NOR2X1 U1043 ( .IN1(n888), .IN2(N270), .OUT(n896) );
  INVX1 U1044 ( .IN(Exc_Ack), .OUT(n889) );
  NOR2X1 U1045 ( .IN1(n1104), .IN2(n889), .OUT(n893) );
  OAI21 U1046 ( .IN1(n222), .IN2(n896), .IN3(n890), .OUT(n1101) );
  AOI22 U1047 ( .IN1(Exc_value[1]), .IN2(n893), .IN3(n242), .IN4(n891), .OUT(
        n892) );
  OAI21 U1048 ( .IN1(n819), .IN2(n1146), .IN3(n892), .OUT(n1093) );
  AOI22 U1049 ( .IN1(n823), .IN2(n894), .IN3(n893), .IN4(Exc_value[0]), .OUT(
        n895) );
  OAI21 U1050 ( .IN1(n896), .IN2(n243), .IN3(n895), .OUT(n1092) );
  OAI21 U1051 ( .IN1(n241), .IN2(n897), .IN3(n285), .OUT(n898) );
  OAI21 U1052 ( .IN1(n898), .IN2(n245), .IN3(n1130), .OUT(n1091) );
  AOI22 U1053 ( .IN1(n821), .IN2(Datain2[0]), .IN3(n822), .IN4(Datain1[0]), 
        .OUT(n899) );
  OAI21 U1054 ( .IN1(n973), .IN2(n219), .IN3(n899), .OUT(n1089) );
  AOI22 U1055 ( .IN1(n821), .IN2(Datain2[1]), .IN3(n822), .IN4(Datain1[1]), 
        .OUT(n900) );
  OAI21 U1056 ( .IN1(n973), .IN2(n218), .IN3(n900), .OUT(n1088) );
  AOI22 U1057 ( .IN1(n821), .IN2(Datain2[2]), .IN3(n822), .IN4(Datain1[2]), 
        .OUT(n901) );
  OAI21 U1058 ( .IN1(n973), .IN2(n217), .IN3(n901), .OUT(n1087) );
  AOI22 U1059 ( .IN1(n821), .IN2(Datain2[3]), .IN3(n822), .IN4(Datain1[3]), 
        .OUT(n902) );
  OAI21 U1060 ( .IN1(n973), .IN2(n216), .IN3(n902), .OUT(n1086) );
  AOI22 U1061 ( .IN1(n821), .IN2(Datain2[4]), .IN3(n822), .IN4(Datain1[4]), 
        .OUT(n903) );
  OAI21 U1062 ( .IN1(n973), .IN2(n215), .IN3(n903), .OUT(n1085) );
  AOI22 U1063 ( .IN1(n821), .IN2(Datain2[5]), .IN3(n822), .IN4(n273), .OUT(
        n904) );
  OAI21 U1064 ( .IN1(n973), .IN2(n214), .IN3(n904), .OUT(n1084) );
  AOI22 U1065 ( .IN1(n821), .IN2(Datain2[6]), .IN3(n822), .IN4(Datain1[6]), 
        .OUT(n905) );
  OAI21 U1066 ( .IN1(n973), .IN2(n213), .IN3(n905), .OUT(n1083) );
  NAND3X1 U1067 ( .IN1(n200), .IN2(n906), .IN3(n199), .OUT(n907) );
  NOR2X1 U1068 ( .IN1(Datain1[9]), .IN2(n907), .OUT(n910) );
  NAND3X1 U1069 ( .IN1(n196), .IN2(n181), .IN3(n194), .OUT(n908) );
  NOR2X1 U1070 ( .IN1(DP_OP_982J1_125_6202_n91), .IN2(n908), .OUT(n909) );
  AOI21 U1071 ( .IN1(n822), .IN2(n944), .IN3(n821), .OUT(n911) );
  OAI21 U1072 ( .IN1(n973), .IN2(n212), .IN3(n911), .OUT(n1082) );
  NOR2X1 U1073 ( .IN1(N423), .IN2(N421), .OUT(n913) );
  NOR2X1 U1074 ( .IN1(N422), .IN2(N424), .OUT(n912) );
  NOR2X1 U1075 ( .IN1(N425), .IN2(n914), .OUT(n999) );
  NAND2X1 U1076 ( .IN1(N420), .IN2(n999), .OUT(n916) );
  NOR2X1 U1077 ( .IN1(n1001), .IN2(n916), .OUT(n977) );
  AOI22 U1078 ( .IN1(N159), .IN2(n273), .IN3(n271), .IN4(n1044), .OUT(n917) );
  NAND3X1 U1079 ( .IN1(Datain1[4]), .IN2(N155), .IN3(N160), .OUT(n942) );
  AOI22 U1080 ( .IN1(n977), .IN2(n1031), .IN3(n250), .IN4(n1052), .OUT(n950)
         );
  NOR2X1 U1081 ( .IN1(DP_OP_982J1_125_6202_n101), .IN2(
        DP_OP_982J1_125_6202_n102), .OUT(n918) );
  NAND3X1 U1082 ( .IN1(n918), .IN2(n179), .IN3(n176), .OUT(n919) );
  NOR2X1 U1083 ( .IN1(Datain2[7]), .IN2(n919), .OUT(n921) );
  NOR2X1 U1084 ( .IN1(DP_OP_982J1_125_6202_n97), .IN2(
        DP_OP_982J1_125_6202_n100), .OUT(n920) );
  NAND3X1 U1085 ( .IN1(n921), .IN2(n920), .IN3(n178), .OUT(n978) );
  NOR2X1 U1086 ( .IN1(n1116), .IN2(n978), .OUT(n983) );
  INVX1 U1087 ( .IN(Datain2[5]), .OUT(n984) );
  NOR2X1 U1088 ( .IN1(n984), .IN2(n270), .OUT(n960) );
  AOI22 U1089 ( .IN1(n270), .IN2(Datain2[6]), .IN3(Datain2[4]), .IN4(N148), 
        .OUT(n1015) );
  AOI22 U1090 ( .IN1(n157), .IN2(n923), .IN3(n1015), .IN4(N143), .OUT(n928) );
  NAND2X1 U1091 ( .IN1(Datain2[4]), .IN2(N148), .OUT(n926) );
  AOI22 U1092 ( .IN1(n157), .IN2(n959), .IN3(n270), .IN4(Datain2[6]), .OUT(
        n925) );
  OAI21 U1093 ( .IN1(n157), .IN2(n926), .IN3(n925), .OUT(n927) );
  AOI22 U1094 ( .IN1(n983), .IN2(n928), .IN3(n1053), .IN4(n927), .OUT(n1027)
         );
  NOR2X1 U1095 ( .IN1(N367), .IN2(N365), .OUT(n930) );
  NOR2X1 U1096 ( .IN1(N366), .IN2(N368), .OUT(n929) );
  NOR2X1 U1097 ( .IN1(n931), .IN2(N369), .OUT(n932) );
  NAND2X1 U1098 ( .IN1(N364), .IN2(n932), .OUT(n958) );
  INVX1 U1099 ( .IN(n932), .OUT(n987) );
  NOR2X1 U1100 ( .IN1(n157), .IN2(n985), .OUT(n975) );
  INVX1 U1101 ( .IN(Datain2[2]), .OUT(n952) );
  INVX1 U1102 ( .IN(Datain2[0]), .OUT(n933) );
  AOI22 U1103 ( .IN1(n270), .IN2(n952), .IN3(n933), .IN4(N148), .OUT(n936) );
  NOR2X1 U1104 ( .IN1(N143), .IN2(n985), .OUT(n1018) );
  INVX1 U1105 ( .IN(Datain2[3]), .OUT(n935) );
  INVX1 U1106 ( .IN(Datain2[1]), .OUT(n934) );
  AOI22 U1107 ( .IN1(n270), .IN2(n935), .IN3(n934), .IN4(N148), .OUT(n954) );
  AOI22 U1108 ( .IN1(n975), .IN2(n936), .IN3(n1018), .IN4(n954), .OUT(n937) );
  OAI21 U1109 ( .IN1(n1027), .IN2(n958), .IN3(n937), .OUT(n940) );
  NOR2X1 U1110 ( .IN1(n998), .IN2(n1001), .OUT(n1038) );
  INVX1 U1111 ( .IN(n1038), .OUT(n951) );
  AOI22 U1112 ( .IN1(Datain1[3]), .IN2(n1019), .IN3(n1045), .IN4(Datain1[1]), 
        .OUT(n956) );
  AOI22 U1113 ( .IN1(n1019), .IN2(Datain1[2]), .IN3(n1045), .IN4(Datain1[0]), 
        .OUT(n938) );
  AOI22 U1114 ( .IN1(N159), .IN2(n956), .IN3(n938), .IN4(N155), .OUT(n939) );
  NOR2X1 U1115 ( .IN1(n940), .IN2(n939), .OUT(n949) );
  NOR2X1 U1116 ( .IN1(N159), .IN2(N420), .OUT(n995) );
  AOI22 U1117 ( .IN1(n271), .IN2(Datain1[2]), .IN3(Datain1[0]), .IN4(N160), 
        .OUT(n941) );
  AOI22 U1118 ( .IN1(n271), .IN2(Datain1[3]), .IN3(Datain1[1]), .IN4(N160), 
        .OUT(n969) );
  NOR2X1 U1119 ( .IN1(N155), .IN2(N420), .OUT(n968) );
  AOI22 U1120 ( .IN1(n995), .IN2(n941), .IN3(n969), .IN4(n968), .OUT(n947) );
  NOR2X1 U1121 ( .IN1(n271), .IN2(N155), .OUT(n1119) );
  NOR2X1 U1122 ( .IN1(N160), .IN2(N159), .OUT(n993) );
  OAI21 U1123 ( .IN1(n964), .IN2(n1011), .IN3(n942), .OUT(n943) );
  AOI21 U1124 ( .IN1(n1119), .IN2(n273), .IN3(n943), .OUT(n1029) );
  NAND3X1 U1125 ( .IN1(n821), .IN2(n999), .IN3(n945), .OUT(n1008) );
  AOI21 U1126 ( .IN1(N420), .IN2(n1029), .IN3(n1008), .OUT(n946) );
  NAND3X1 U1127 ( .IN1(n950), .IN2(n949), .IN3(n948), .OUT(n1080) );
  AOI22 U1128 ( .IN1(n271), .IN2(Datain1[4]), .IN3(Datain1[2]), .IN4(N160), 
        .OUT(n967) );
  NOR2X1 U1129 ( .IN1(n951), .IN2(n967), .OUT(n980) );
  INVX1 U1130 ( .IN(Datain2[4]), .OUT(n953) );
  AOI22 U1131 ( .IN1(n270), .IN2(n953), .IN3(n952), .IN4(N148), .OUT(n974) );
  AOI22 U1132 ( .IN1(n975), .IN2(n954), .IN3(n1018), .IN4(n974), .OUT(n955) );
  OAI21 U1133 ( .IN1(n956), .IN2(N159), .IN3(n955), .OUT(n957) );
  NAND3X1 U1134 ( .IN1(n822), .IN2(Datain2[6]), .IN3(N148), .OUT(n962) );
  AOI22 U1135 ( .IN1(n983), .IN2(n960), .IN3(n1053), .IN4(n959), .OUT(n961) );
  AOI22 U1136 ( .IN1(n157), .IN2(n962), .IN3(n961), .IN4(N143), .OUT(n1034) );
  NAND2X1 U1137 ( .IN1(n1119), .IN2(Datain1[6]), .OUT(n963) );
  NAND3X1 U1138 ( .IN1(n964), .IN2(n965), .IN3(n963), .OUT(n1037) );
  AOI22 U1139 ( .IN1(Datain1[6]), .IN2(n1119), .IN3(n966), .IN4(N160), .OUT(
        n1035) );
  AOI22 U1140 ( .IN1(N420), .IN2(n1035), .IN3(n968), .IN4(n967), .OUT(n971) );
  AOI21 U1141 ( .IN1(n995), .IN2(n969), .IN3(n1008), .OUT(n970) );
  AOI22 U1142 ( .IN1(n977), .IN2(n1037), .IN3(n971), .IN4(n970), .OUT(n972) );
  NOR2X1 U1143 ( .IN1(n271), .IN2(n1011), .OUT(n976) );
  AOI22 U1144 ( .IN1(n977), .IN2(n976), .IN3(n975), .IN4(n974), .OUT(n1007) );
  OAI21 U1145 ( .IN1(N143), .IN2(n978), .IN3(n822), .OUT(n1041) );
  NAND2X1 U1146 ( .IN1(Datain2[6]), .IN2(N148), .OUT(n979) );
  NOR2X1 U1147 ( .IN1(n1041), .IN2(n979), .OUT(n982) );
  AOI22 U1148 ( .IN1(n982), .IN2(n981), .IN3(n980), .IN4(N155), .OUT(n1006) );
  NAND2X1 U1149 ( .IN1(Datain2[3]), .IN2(n983), .OUT(n992) );
  NOR2X1 U1150 ( .IN1(n985), .IN2(n984), .OUT(n989) );
  OAI21 U1151 ( .IN1(N364), .IN2(Datain2[3]), .IN3(n1053), .OUT(n986) );
  NOR2X1 U1152 ( .IN1(n987), .IN2(n986), .OUT(n988) );
  AOI22 U1153 ( .IN1(n270), .IN2(n989), .IN3(n988), .IN4(N148), .OUT(n990) );
  OAI21 U1154 ( .IN1(n1051), .IN2(n992), .IN3(n990), .OUT(n1021) );
  NOR2X1 U1155 ( .IN1(n271), .IN2(Datain1[2]), .OUT(n994) );
  INVX1 U1156 ( .IN(Datain1[4]), .OUT(n1012) );
  AOI22 U1157 ( .IN1(n995), .IN2(n994), .IN3(n993), .IN4(n1012), .OUT(n997) );
  AOI22 U1158 ( .IN1(n271), .IN2(n273), .IN3(Datain1[3]), .IN4(N160), .OUT(
        n1010) );
  NAND3X1 U1159 ( .IN1(Datain1[6]), .IN2(N155), .IN3(N160), .OUT(n1046) );
  AOI22 U1160 ( .IN1(N159), .IN2(n1010), .IN3(N420), .IN4(n1046), .OUT(n996)
         );
  OAI21 U1161 ( .IN1(Datain1[3]), .IN2(N420), .IN3(n999), .OUT(n1000) );
  AOI22 U1162 ( .IN1(N159), .IN2(n1016), .IN3(n1052), .IN4(n249), .OUT(n1002)
         );
  OAI21 U1163 ( .IN1(n1008), .IN2(n1003), .IN3(n1002), .OUT(n1004) );
  AOI21 U1164 ( .IN1(n157), .IN2(n1021), .IN3(n1004), .OUT(n1005) );
  NAND3X1 U1165 ( .IN1(n1005), .IN2(n1006), .IN3(n1007), .OUT(n1078) );
  NOR2X1 U1166 ( .IN1(n1008), .IN2(N420), .OUT(n1048) );
  INVX1 U1167 ( .IN(n1048), .OUT(n1009) );
  AOI21 U1168 ( .IN1(n1010), .IN2(N155), .IN3(n1009), .OUT(n1014) );
  NOR2X1 U1169 ( .IN1(N155), .IN2(N160), .OUT(n1109) );
  AOI22 U1170 ( .IN1(n1119), .IN2(n1012), .IN3(n1109), .IN4(n1011), .OUT(n1013) );
  AOI22 U1171 ( .IN1(n1014), .IN2(n1013), .IN3(n1052), .IN4(n221), .OUT(n1026)
         );
  AOI22 U1172 ( .IN1(n1018), .IN2(n1017), .IN3(n1016), .IN4(N155), .OUT(n1025)
         );
  AOI22 U1173 ( .IN1(n1019), .IN2(Datain1[6]), .IN3(n1045), .IN4(Datain1[4]), 
        .OUT(n1020) );
  AOI22 U1174 ( .IN1(N159), .IN2(n1022), .IN3(N143), .IN4(n1021), .OUT(n1023)
         );
  NAND3X1 U1175 ( .IN1(n1026), .IN2(n1025), .IN3(n1023), .OUT(n1077) );
  INVX1 U1176 ( .IN(n1027), .OUT(n1028) );
  AOI22 U1177 ( .IN1(n1112), .IN2(n1028), .IN3(n1052), .IN4(n248), .OUT(n1033)
         );
  AOI22 U1178 ( .IN1(n1038), .IN2(n1031), .IN3(n1048), .IN4(n1030), .OUT(n1032) );
  AOI22 U1179 ( .IN1(n1034), .IN2(n1112), .IN3(n1052), .IN4(n224), .OUT(n1040)
         );
  AOI22 U1180 ( .IN1(n1038), .IN2(n1037), .IN3(n1048), .IN4(n1036), .OUT(n1039) );
  INVX1 U1181 ( .IN(Datain2[6]), .OUT(n1042) );
  AOI21 U1182 ( .IN1(N143), .IN2(n1042), .IN3(n1041), .OUT(n1043) );
  AOI22 U1183 ( .IN1(n1045), .IN2(n1044), .IN3(n1117), .IN4(n1043), .OUT(n1050) );
  AOI22 U1184 ( .IN1(n1048), .IN2(n1047), .IN3(n1052), .IN4(n247), .OUT(n1049)
         );
  NOR2X1 U1185 ( .IN1(n157), .IN2(n1051), .OUT(n1056) );
  AOI22 U1186 ( .IN1(n1056), .IN2(n1053), .IN3(Op2_Mantissa_reg_7_), .IN4(
        n1052), .OUT(n1054) );
  OAI21 U1187 ( .IN1(N159), .IN2(n1055), .IN3(n1054), .OUT(n1073) );
  NOR2X1 U1188 ( .IN1(n1056), .IN2(n1116), .OUT(n1057) );
  AOI22 U1189 ( .IN1(n821), .IN2(N430), .IN3(N376), .IN4(n1057), .OUT(n1108)
         );
  NOR2X1 U1190 ( .IN1(n211), .IN2(n240), .OUT(n1128) );
  MUX2X1 U1191 ( .IN1(add_x_35_A_2_), .IN2(n226), .S(n1128), .OUT(n1106) );
  OAI21 U1192 ( .IN1(n1145), .IN2(n1059), .IN3(n285), .OUT(n1105) );
  NAND2X1 U1193 ( .IN1(n1108), .IN2(n1107), .OUT(n1072) );
  AOI21 U1194 ( .IN1(n1120), .IN2(n1110), .IN3(n1118), .OUT(n1114) );
  AOI21 U1195 ( .IN1(n1112), .IN2(n1111), .IN3(n1116), .OUT(n1113) );
  AOI22 U1196 ( .IN1(N445), .IN2(n1114), .IN3(N392), .IN4(n1113), .OUT(n1115)
         );
  NOR2X1 U1197 ( .IN1(n1117), .IN2(n1116), .OUT(n1122) );
  AOI21 U1198 ( .IN1(n1120), .IN2(n1119), .IN3(n1118), .OUT(n1121) );
  AOI22 U1199 ( .IN1(N384), .IN2(n1122), .IN3(N437), .IN4(n1121), .OUT(n1124)
         );
  NAND2X1 U1200 ( .IN1(n1124), .IN2(n1123), .OUT(n1070) );
  OAI21 U1201 ( .IN1(n1146), .IN2(n1127), .IN3(n1126), .OUT(n1060) );
  NOR2X1 U1202 ( .IN1(n250), .IN2(n1137), .OUT(n1136) );
  NAND2X1 U1203 ( .IN1(add_x_35_A_4_), .IN2(n1136), .OUT(n1135) );
  NOR2X1 U1204 ( .IN1(n249), .IN2(n1135), .OUT(n1134) );
  NOR2X1 U1205 ( .IN1(n248), .IN2(n1133), .OUT(n1132) );
  NOR2X1 U1206 ( .IN1(n247), .IN2(n1131), .OUT(n1129) );
  AOI22 U1207 ( .IN1(n823), .IN2(n1140), .IN3(Debug_reg[2]), .IN4(n1144), 
        .OUT(n1141) );
  AOI22 U1208 ( .IN1(n823), .IN2(n1142), .IN3(Debug_reg[1]), .IN4(n1144), 
        .OUT(n1143) );
  OAI21 U1209 ( .IN1(n1147), .IN2(n246), .IN3(n1146), .OUT(n103) );
  MUX2X1 U1210 ( .IN1(n1168), .IN2(n1169), .S(N144), .OUT(n1148) );
  MUX2X1 U1211 ( .IN1(n1170), .IN2(n1171), .S(N144), .OUT(n1149) );
  MUX2X1 U1212 ( .IN1(n1172), .IN2(n1173), .S(N144), .OUT(n1150) );
  MUX2X1 U1213 ( .IN1(n1174), .IN2(n1175), .S(N144), .OUT(n1151) );
  MUX2X1 U1214 ( .IN1(n1148), .IN2(n1149), .S(N145), .OUT(n1152) );
  MUX2X1 U1215 ( .IN1(n1152), .IN2(n1153), .S(N146), .OUT(N376) );
  MUX2X1 U1216 ( .IN1(Datain2[0]), .IN2(Datain2[1]), .S(n157), .OUT(n1154) );
  MUX2X1 U1217 ( .IN1(Datain2[2]), .IN2(Datain2[3]), .S(n157), .OUT(n1155) );
  MUX2X1 U1218 ( .IN1(Datain2[4]), .IN2(Datain2[5]), .S(N147), .OUT(n1156) );
  MUX2X1 U1219 ( .IN1(Datain2[6]), .IN2(Datain2[7]), .S(N147), .OUT(n1157) );
  MUX2X1 U1220 ( .IN1(Datain2[8]), .IN2(DP_OP_982J1_125_6202_n97), .S(N147), 
        .OUT(n1158) );
  MUX2X1 U1221 ( .IN1(Datain2[10]), .IN2(Datain2[11]), .S(N147), .OUT(n1159)
         );
  MUX2X1 U1222 ( .IN1(DP_OP_982J1_125_6202_n100), .IN2(
        DP_OP_982J1_125_6202_n101), .S(n157), .OUT(n1160) );
  MUX2X1 U1223 ( .IN1(DP_OP_982J1_125_6202_n102), .IN2(Datain2[15]), .S(n157), 
        .OUT(n1161) );
  MUX2X1 U1224 ( .IN1(n1154), .IN2(n1155), .S(N148), .OUT(n1162) );
  MUX2X1 U1225 ( .IN1(n1156), .IN2(n1157), .S(N148), .OUT(n1163) );
  MUX2X1 U1226 ( .IN1(n1158), .IN2(n1159), .S(N148), .OUT(n1164) );
  MUX2X1 U1227 ( .IN1(n1160), .IN2(n1161), .S(N148), .OUT(n1165) );
  MUX2X1 U1228 ( .IN1(n1162), .IN2(n1163), .S(N149), .OUT(n1166) );
  MUX2X1 U1229 ( .IN1(n1166), .IN2(n1167), .S(N150), .OUT(N384) );
  MUX2X1 U1230 ( .IN1(Datain2[0]), .IN2(Datain2[1]), .S(N143), .OUT(n1168) );
  MUX2X1 U1231 ( .IN1(Datain2[2]), .IN2(Datain2[3]), .S(N143), .OUT(n1169) );
  MUX2X1 U1232 ( .IN1(Datain2[4]), .IN2(Datain2[5]), .S(N143), .OUT(n1170) );
  MUX2X1 U1233 ( .IN1(Datain2[6]), .IN2(Datain2[7]), .S(N143), .OUT(n1171) );
  MUX2X1 U1234 ( .IN1(Datain2[8]), .IN2(DP_OP_982J1_125_6202_n97), .S(N143), 
        .OUT(n1172) );
  MUX2X1 U1235 ( .IN1(Datain2[10]), .IN2(Datain2[11]), .S(N143), .OUT(n1173)
         );
  MUX2X1 U1236 ( .IN1(DP_OP_982J1_125_6202_n100), .IN2(
        DP_OP_982J1_125_6202_n101), .S(N143), .OUT(n1174) );
  MUX2X1 U1237 ( .IN1(DP_OP_982J1_125_6202_n102), .IN2(Datain2[15]), .S(N143), 
        .OUT(n1175) );
  MUX2X1 U1238 ( .IN1(n1168), .IN2(n1169), .S(N152), .OUT(n1176) );
  MUX2X1 U1239 ( .IN1(n1170), .IN2(n1171), .S(N152), .OUT(n1177) );
  MUX2X1 U1240 ( .IN1(n1172), .IN2(n1173), .S(N152), .OUT(n1178) );
  MUX2X1 U1241 ( .IN1(n1174), .IN2(n1175), .S(N152), .OUT(n1179) );
  MUX2X1 U1242 ( .IN1(n1176), .IN2(n1177), .S(N153), .OUT(n1180) );
  MUX2X1 U1243 ( .IN1(n1180), .IN2(n1181), .S(N154), .OUT(N392) );
  MUX2X1 U1244 ( .IN1(n1190), .IN2(n1191), .S(N156), .OUT(n1182) );
  MUX2X1 U1245 ( .IN1(n1192), .IN2(n1193), .S(N156), .OUT(n1183) );
  MUX2X1 U1246 ( .IN1(n1194), .IN2(n1195), .S(N156), .OUT(n1184) );
  MUX2X1 U1247 ( .IN1(n1196), .IN2(n1197), .S(N156), .OUT(n1185) );
  MUX2X1 U1248 ( .IN1(n1182), .IN2(n1183), .S(N157), .OUT(n1186) );
  MUX2X1 U1249 ( .IN1(n1184), .IN2(n1185), .S(N157), .OUT(n1187) );
  MUX2X1 U1250 ( .IN1(n1186), .IN2(n1187), .S(N158), .OUT(N430) );
  MUX2X1 U1251 ( .IN1(n1188), .IN2(n1189), .S(N162), .OUT(N437) );
  MUX2X1 U1252 ( .IN1(Datain1[0]), .IN2(Datain1[1]), .S(N155), .OUT(n1190) );
  MUX2X1 U1253 ( .IN1(Datain1[2]), .IN2(Datain1[3]), .S(N155), .OUT(n1191) );
  MUX2X1 U1254 ( .IN1(Datain1[4]), .IN2(n273), .S(N155), .OUT(n1192) );
  MUX2X1 U1255 ( .IN1(Datain1[6]), .IN2(Datain1[7]), .S(N155), .OUT(n1193) );
  MUX2X1 U1256 ( .IN1(Datain1[8]), .IN2(Datain1[9]), .S(N155), .OUT(n1194) );
  MUX2X1 U1257 ( .IN1(Datain1[10]), .IN2(DP_OP_982J1_125_6202_n91), .S(N155), 
        .OUT(n1195) );
  MUX2X1 U1258 ( .IN1(Datain1[12]), .IN2(Datain1[13]), .S(N155), .OUT(n1196)
         );
  MUX2X1 U1259 ( .IN1(Datain1[14]), .IN2(Datain1[15]), .S(N155), .OUT(n1197)
         );
  MUX2X1 U1260 ( .IN1(n1190), .IN2(n1191), .S(N164), .OUT(n1198) );
  MUX2X1 U1261 ( .IN1(n1192), .IN2(n1193), .S(N164), .OUT(n1199) );
  MUX2X1 U1262 ( .IN1(n1194), .IN2(n1195), .S(N164), .OUT(n1200) );
  MUX2X1 U1263 ( .IN1(n1196), .IN2(n1197), .S(N164), .OUT(n1201) );
  MUX2X1 U1264 ( .IN1(n1198), .IN2(n1199), .S(N165), .OUT(n1202) );
  MUX2X1 U1265 ( .IN1(n1200), .IN2(n1201), .S(N165), .OUT(n1203) );
  MUX2X1 U1266 ( .IN1(n1202), .IN2(n1203), .S(N166), .OUT(N445) );
endmodule


module Mul_cntrl ( CLK, Datain1, Datain2, Data_valid, Dataout, Dataout_valid, 
        Exc, Mode, Debug, Multi_datain1, Multi_datain2, Multi_dataout, 
        Multi_ack, ExcCheck_valid, ExcCheck_Datain, Exc_value, RSTn_BAR, 
        Multi_valid_BAR, Exc_Ack_BAR );
  input [15:0] Datain1;
  input [15:0] Datain2;
  output [15:0] Dataout;
  output [2:0] Exc;
  input [2:0] Mode;
  output [4:0] Debug;
  output [7:0] Multi_datain1;
  output [7:0] Multi_datain2;
  input [15:0] Multi_dataout;
  output [15:0] ExcCheck_Datain;
  input [2:0] Exc_value;
  input CLK, Data_valid, Multi_ack, RSTn_BAR, Exc_Ack_BAR;
  output Dataout_valid, ExcCheck_valid, Multi_valid_BAR;
  wire   Debug_valid_reg, Final_Sign_reg, G_reg, T_reg, N89, N90, N384, N385,
         N386, N387, N388, N389, N390, N391, N392, C276_DATA3_0, C276_DATA3_1,
         C276_DATA3_2, C276_DATA3_3, C276_DATA3_5, C276_DATA3_6, C276_DATA3_7,
         n64, n94, n96, n124, n125, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n144, n145, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n213, n214, n215, n667, n703, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, C1_Z_3,
         C1_Z_2, C1_Z_1, C1_Z_0, RSOP_428_C1_Z_0, DP_OP_433_158_7755_n75,
         DP_OP_433_158_7755_n74, DP_OP_433_158_7755_n73,
         DP_OP_433_158_7755_n69, DP_OP_433_158_7755_n68,
         DP_OP_433_158_7755_n67, DP_OP_433_158_7755_n66,
         DP_OP_433_158_7755_n65, DP_OP_433_158_7755_n64,
         DP_OP_433_158_7755_n63, DP_OP_433_158_7755_n62,
         DP_OP_433_158_7755_n61, DP_OP_433_158_7755_n60,
         DP_OP_433_158_7755_n59, DP_OP_433_158_7755_n58,
         DP_OP_433_158_7755_n57, DP_OP_433_158_7755_n56,
         DP_OP_433_158_7755_n52, DP_OP_433_158_7755_n48,
         DP_OP_433_158_7755_n46, DP_OP_433_158_7755_n43,
         DP_OP_433_158_7755_n42, DP_OP_433_158_7755_n38,
         DP_OP_433_158_7755_n37, DP_OP_433_158_7755_n33,
         DP_OP_433_158_7755_n19, DP_OP_433_158_7755_n18,
         DP_OP_433_158_7755_n17, DP_OP_433_158_7755_n16,
         DP_OP_433_158_7755_n13, DP_OP_433_158_7755_n10, DP_OP_433_158_7755_n7,
         DP_OP_433_158_7755_n1, DP_OP_357J3_124_4634_n66,
         DP_OP_357J3_124_4634_n65, DP_OP_357J3_124_4634_n58,
         DP_OP_357J3_124_4634_n29, DP_OP_357J3_124_4634_n28,
         DP_OP_357J3_124_4634_n27, DP_OP_357J3_124_4634_n26,
         DP_OP_357J3_124_4634_n25, DP_OP_357J3_124_4634_n24,
         DP_OP_357J3_124_4634_n23, DP_OP_357J3_124_4634_n22,
         DP_OP_357J3_124_4634_n21, DP_OP_357J3_124_4634_n20,
         DP_OP_357J3_124_4634_n19, DP_OP_357J3_124_4634_n18,
         DP_OP_357J3_124_4634_n17, DP_OP_357J3_124_4634_n15,
         DP_OP_357J3_124_4634_n13, DP_OP_357J3_124_4634_n12,
         DP_OP_357J3_124_4634_n11, DP_OP_357J3_124_4634_n10,
         DP_OP_357J3_124_4634_n9, DP_OP_357J3_124_4634_n8,
         DP_OP_357J3_124_4634_n7, DP_OP_357J3_124_4634_n6,
         DP_OP_357J3_124_4634_n5, DP_OP_357J3_124_4634_n4, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n95, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n122, n123, n126, n127, n143, n146, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940;
  wire   [2:0] StateMC;
  wire   [3:0] Debug_reg;
  wire   [8:0] Final_Exponent_reg;
  wire   [7:0] Op1_Mantissa_reg;
  wire   [7:0] Op2_Mantissa_reg;
  wire   [6:0] Final_Mantissa_reg;

  DFFRX1 T_reg_reg ( .D(n124), .CLK(CLK), .CLRB(n64), .Q(T_reg), .QB(n114) );
  DFFRX1 exc_reg_reg_2_ ( .D(n667), .CLK(CLK), .CLRB(n64), .Q(n213), .QB(n108)
         );
  DFFRX1 StateMC_reg_0_ ( .D(n703), .CLK(CLK), .CLRB(n64), .Q(n104), .QB(
        StateMC[0]) );
  DFFRX1 StateMC_reg_1_ ( .D(N89), .CLK(CLK), .CLRB(n64), .Q(StateMC[1]), .QB(
        n105) );
  DFFRX1 StateMC_reg_2_ ( .D(N90), .CLK(CLK), .CLRB(n64), .Q(StateMC[2]), .QB(
        n99) );
  DFFRX1 Op1_Mantissa_reg_reg_0_ ( .D(n147), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[0]) );
  DFFRX1 Op1_Mantissa_reg_reg_1_ ( .D(n148), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[1]) );
  DFFRX1 Op1_Mantissa_reg_reg_2_ ( .D(n149), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[2]) );
  DFFRX1 Op1_Mantissa_reg_reg_3_ ( .D(n150), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[3]) );
  DFFRX1 Op1_Mantissa_reg_reg_4_ ( .D(n151), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[4]) );
  DFFRX1 Op1_Mantissa_reg_reg_5_ ( .D(n152), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[5]) );
  DFFRX1 Op1_Mantissa_reg_reg_6_ ( .D(n153), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[6]) );
  DFFRX1 Op1_Mantissa_reg_reg_7_ ( .D(n154), .CLK(CLK), .CLRB(n64), .Q(
        Op1_Mantissa_reg[7]) );
  DFFRX1 Op2_Mantissa_reg_reg_0_ ( .D(n155), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[0]) );
  DFFRX1 Op2_Mantissa_reg_reg_1_ ( .D(n156), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[1]) );
  DFFRX1 Op2_Mantissa_reg_reg_2_ ( .D(n157), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[2]) );
  DFFRX1 Op2_Mantissa_reg_reg_3_ ( .D(n158), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[3]) );
  DFFRX1 Op2_Mantissa_reg_reg_4_ ( .D(n159), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[4]) );
  DFFRX1 Op2_Mantissa_reg_reg_5_ ( .D(n160), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[5]) );
  DFFRX1 Op2_Mantissa_reg_reg_6_ ( .D(n161), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[6]) );
  DFFRX1 Op2_Mantissa_reg_reg_7_ ( .D(n881), .CLK(CLK), .CLRB(n64), .Q(
        Op2_Mantissa_reg[7]) );
  DFFRX1 exc_reg_reg_0_ ( .D(n882), .CLK(CLK), .CLRB(n64), .QB(n215) );
  DFFRX1 Final_Exponent_reg_reg_8_ ( .D(n94), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[8]), .QB(n119) );
  DFFRX1 exc_reg_reg_1_ ( .D(n883), .CLK(CLK), .CLRB(n64), .Q(n120), .QB(n214)
         );
  DFFRX1 Final_Exponent_reg_reg_7_ ( .D(n872), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[7]), .QB(n117) );
  DFFRX1 Final_Exponent_reg_reg_6_ ( .D(n873), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[6]), .QB(n100) );
  DFFRX1 Final_Exponent_reg_reg_5_ ( .D(n874), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[5]), .QB(n116) );
  DFFRX1 Final_Exponent_reg_reg_4_ ( .D(n875), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[4]), .QB(n118) );
  DFFRX1 Final_Exponent_reg_reg_3_ ( .D(n876), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[3]), .QB(n102) );
  DFFRX1 Final_Exponent_reg_reg_2_ ( .D(n877), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[2]), .QB(n98) );
  DFFRX1 Final_Exponent_reg_reg_1_ ( .D(n878), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[1]), .QB(n97) );
  DFFRX1 Final_Exponent_reg_reg_0_ ( .D(n879), .CLK(CLK), .CLRB(n64), .Q(
        Final_Exponent_reg[0]), .QB(n103) );
  DFFRX1 Debug_valid_reg_reg ( .D(n96), .CLK(CLK), .CLRB(n64), .Q(
        Debug_valid_reg) );
  DFFRX1 Final_Mantissa_reg_reg_0_ ( .D(n871), .CLK(CLK), .CLRB(n64), .Q(
        Final_Mantissa_reg[0]), .QB(n107) );
  DFFRX1 Final_Mantissa_reg_reg_1_ ( .D(n870), .CLK(CLK), .CLRB(n64), .Q(
        Final_Mantissa_reg[1]), .QB(n111) );
  DFFRX1 Final_Mantissa_reg_reg_2_ ( .D(n869), .CLK(CLK), .CLRB(n64), .Q(
        Final_Mantissa_reg[2]), .QB(n109) );
  DFFRX1 Final_Mantissa_reg_reg_3_ ( .D(n868), .CLK(CLK), .CLRB(n64), .Q(
        Final_Mantissa_reg[3]), .QB(n106) );
  DFFRX1 Final_Mantissa_reg_reg_4_ ( .D(n867), .CLK(CLK), .CLRB(n64), .Q(
        Final_Mantissa_reg[4]), .QB(n112) );
  DFFRX1 Final_Mantissa_reg_reg_5_ ( .D(n866), .CLK(CLK), .CLRB(n64), .Q(
        Final_Mantissa_reg[5]), .QB(n110) );
  DFFRX1 Final_Mantissa_reg_reg_6_ ( .D(n865), .CLK(CLK), .CLRB(n64), .Q(
        Final_Mantissa_reg[6]), .QB(n113) );
  DFFRX1 Final_Sign_reg_reg ( .D(n880), .CLK(CLK), .CLRB(n64), .Q(
        Final_Sign_reg) );
  DFFRX1 G_reg_reg ( .D(n125), .CLK(CLK), .CLRB(n64), .Q(G_reg), .QB(n101) );
  DFFRX1 Multi_datain1_reg_7_ ( .D(n163), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[7]) );
  DFFRX1 Multi_datain1_reg_6_ ( .D(n162), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[6]) );
  DFFRX1 Multi_datain1_reg_5_ ( .D(n133), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[5]) );
  DFFRX1 Multi_datain1_reg_4_ ( .D(n132), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[4]) );
  DFFRX1 Multi_datain1_reg_3_ ( .D(n131), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[3]) );
  DFFRX1 Multi_datain1_reg_2_ ( .D(n130), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[2]) );
  DFFRX1 Multi_datain1_reg_1_ ( .D(n129), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[1]) );
  DFFRX1 Multi_datain1_reg_0_ ( .D(n128), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain1[0]) );
  DFFRX1 Multi_datain2_reg_7_ ( .D(n141), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[7]) );
  DFFRX1 Multi_datain2_reg_6_ ( .D(n140), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[6]) );
  DFFRX1 Multi_datain2_reg_5_ ( .D(n139), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[5]) );
  DFFRX1 Multi_datain2_reg_4_ ( .D(n138), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[4]) );
  DFFRX1 Multi_datain2_reg_3_ ( .D(n137), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[3]) );
  DFFRX1 Multi_datain2_reg_2_ ( .D(n136), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[2]) );
  DFFRX1 Multi_datain2_reg_1_ ( .D(n135), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[1]) );
  DFFRX1 Multi_datain2_reg_0_ ( .D(n134), .CLK(CLK), .CLRB(n64), .Q(
        Multi_datain2[0]) );
  DFFRX1 Multi_valid_reg ( .D(n142), .CLK(CLK), .CLRB(n64), .QB(
        Multi_valid_BAR) );
  DFFRX1 ExcCheck_valid_reg ( .D(n864), .CLK(CLK), .CLRB(n64), .Q(
        ExcCheck_valid) );
  DFFRX1 Debug_reg_reg_3_ ( .D(n145), .CLK(CLK), .CLRB(n64), .Q(Debug_reg[3])
         );
  DFFRX1 Debug_reg_reg_2_ ( .D(n144), .CLK(CLK), .CLRB(n64), .Q(Debug_reg[2])
         );
  DFFRX1 Debug_reg_reg_1_ ( .D(n862), .CLK(CLK), .CLRB(n64), .Q(Debug_reg[1])
         );
  DFFRX1 Debug_reg_reg_0_ ( .D(n863), .CLK(CLK), .CLRB(n64), .Q(Debug_reg[0]), 
        .QB(n115) );
  NOR2X1 DP_OP_433_158_7755_U80 ( .IN1(Final_Exponent_reg[0]), .IN2(
        DP_OP_433_158_7755_n75), .OUT(DP_OP_433_158_7755_n68) );
  NOR2X1 DP_OP_433_158_7755_U74 ( .IN1(Final_Exponent_reg[1]), .IN2(
        DP_OP_433_158_7755_n74), .OUT(DP_OP_433_158_7755_n66) );
  OAI21 DP_OP_433_158_7755_U71 ( .IN1(DP_OP_433_158_7755_n68), .IN2(
        DP_OP_433_158_7755_n66), .IN3(DP_OP_433_158_7755_n67), .OUT(
        DP_OP_433_158_7755_n65) );
  NOR2X1 DP_OP_433_158_7755_U64 ( .IN1(n204), .IN2(DP_OP_433_158_7755_n73), 
        .OUT(DP_OP_433_158_7755_n62) );
  OAI21 DP_OP_433_158_7755_U61 ( .IN1(DP_OP_433_158_7755_n62), .IN2(
        DP_OP_433_158_7755_n64), .IN3(DP_OP_433_158_7755_n63), .OUT(
        DP_OP_433_158_7755_n61) );
  NOR2X1 DP_OP_433_158_7755_U55 ( .IN1(Final_Exponent_reg[3]), .IN2(n199), 
        .OUT(DP_OP_433_158_7755_n59) );
  OAI21 DP_OP_433_158_7755_U52 ( .IN1(DP_OP_433_158_7755_n63), .IN2(
        DP_OP_433_158_7755_n59), .IN3(DP_OP_433_158_7755_n60), .OUT(
        DP_OP_433_158_7755_n58) );
  NOR2X1 DP_OP_433_158_7755_U51 ( .IN1(DP_OP_433_158_7755_n59), .IN2(
        DP_OP_433_158_7755_n62), .OUT(DP_OP_433_158_7755_n57) );
  AOI21 DP_OP_433_158_7755_U50 ( .IN1(DP_OP_433_158_7755_n57), .IN2(
        DP_OP_433_158_7755_n65), .IN3(DP_OP_433_158_7755_n58), .OUT(
        DP_OP_433_158_7755_n56) );
  NOR2X1 DP_OP_433_158_7755_U49 ( .IN1(DP_OP_433_158_7755_n61), .IN2(
        DP_OP_433_158_7755_n33), .OUT(DP_OP_433_158_7755_n19) );
  NOR2X1 DP_OP_433_158_7755_U48 ( .IN1(DP_OP_433_158_7755_n61), .IN2(
        DP_OP_433_158_7755_n19), .OUT(DP_OP_433_158_7755_n18) );
  NOR2X1 DP_OP_433_158_7755_U47 ( .IN1(DP_OP_433_158_7755_n33), .IN2(
        DP_OP_433_158_7755_n19), .OUT(DP_OP_433_158_7755_n17) );
  NOR2X1 DP_OP_433_158_7755_U46 ( .IN1(DP_OP_433_158_7755_n18), .IN2(
        DP_OP_433_158_7755_n17), .OUT(C276_DATA3_3) );
  NAND2X1 DP_OP_433_158_7755_U41 ( .IN1(DP_OP_433_158_7755_n1), .IN2(n118), 
        .OUT(DP_OP_433_158_7755_n52) );
  NOR2X1 DP_OP_433_158_7755_U29 ( .IN1(DP_OP_433_158_7755_n52), .IN2(
        Final_Exponent_reg[5]), .OUT(DP_OP_433_158_7755_n13) );
  NOR2X1 DP_OP_433_158_7755_U22 ( .IN1(Final_Exponent_reg[6]), .IN2(
        DP_OP_433_158_7755_n48), .OUT(DP_OP_433_158_7755_n43) );
  NOR2X1 DP_OP_433_158_7755_U20 ( .IN1(DP_OP_433_158_7755_n46), .IN2(
        Final_Exponent_reg[6]), .OUT(DP_OP_433_158_7755_n10) );
  NAND2X1 DP_OP_433_158_7755_U12 ( .IN1(n228), .IN2(n227), .OUT(
        DP_OP_433_158_7755_n38) );
  NOR2X1 DP_OP_433_158_7755_U9 ( .IN1(DP_OP_433_158_7755_n42), .IN2(
        Final_Exponent_reg[7]), .OUT(DP_OP_433_158_7755_n7) );
  INVX1 DP_OP_433_158_7755_U32 ( .IN(n227), .OUT(DP_OP_433_158_7755_n48) );
  INVX4 DP_OP_433_158_7755_U82 ( .IN(C1_Z_2), .OUT(DP_OP_433_158_7755_n73) );
  INVX4 DP_OP_433_158_7755_U84 ( .IN(C1_Z_0), .OUT(DP_OP_433_158_7755_n75) );
  INVX4 DP_OP_433_158_7755_U83 ( .IN(C1_Z_1), .OUT(DP_OP_433_158_7755_n74) );
  NANDX2 DP_OP_433_158_7755_U75 ( .IN1(DP_OP_433_158_7755_n74), .IN2(
        Final_Exponent_reg[1]), .OUT(DP_OP_433_158_7755_n67) );
  NANDX2 DP_OP_433_158_7755_U65 ( .IN1(DP_OP_433_158_7755_n73), .IN2(n204), 
        .OUT(DP_OP_433_158_7755_n63) );
  NANDX2 DP_OP_433_158_7755_U56 ( .IN1(n199), .IN2(Final_Exponent_reg[3]), 
        .OUT(DP_OP_433_158_7755_n60) );
  NANDX2 DP_OP_433_158_7755_U40 ( .IN1(DP_OP_433_158_7755_n1), .IN2(
        Final_Exponent_reg[4]), .OUT(DP_OP_433_158_7755_n16) );
  NAND2X1 DP_OP_433_158_7755_U21 ( .IN1(DP_OP_433_158_7755_n1), .IN2(
        DP_OP_433_158_7755_n43), .OUT(DP_OP_433_158_7755_n42) );
  INVX1 DP_OP_433_158_7755_U70 ( .IN(DP_OP_433_158_7755_n65), .OUT(
        DP_OP_433_158_7755_n64) );
  NOR2X1 DP_OP_357J3_124_4634_U18 ( .IN1(Datain2[14]), .IN2(Datain1[14]), 
        .OUT(DP_OP_357J3_124_4634_n15) );
  NOR2X1 DP_OP_357J3_124_4634_U15 ( .IN1(Datain1[14]), .IN2(
        DP_OP_357J3_124_4634_n15), .OUT(DP_OP_357J3_124_4634_n13) );
  NOR2X1 DP_OP_357J3_124_4634_U14 ( .IN1(Datain2[14]), .IN2(
        DP_OP_357J3_124_4634_n15), .OUT(DP_OP_357J3_124_4634_n12) );
  NOR2X1 DP_OP_357J3_124_4634_U13 ( .IN1(DP_OP_357J3_124_4634_n13), .IN2(
        DP_OP_357J3_124_4634_n12), .OUT(DP_OP_357J3_124_4634_n17) );
  FULLADD DP_OP_357J3_124_4634_U12 ( .A(DP_OP_357J3_124_4634_n65), .B(
        Datain2[7]), .CIN(RSOP_428_C1_Z_0), .COUT(DP_OP_357J3_124_4634_n11), 
        .SUM(N384) );
  FULLADD DP_OP_357J3_124_4634_U11 ( .A(n69), .B(n65), .CIN(
        DP_OP_357J3_124_4634_n29), .COUT(DP_OP_357J3_124_4634_n10), .SUM(N385)
         );
  FULLADD DP_OP_357J3_124_4634_U10 ( .A(DP_OP_357J3_124_4634_n27), .B(
        DP_OP_357J3_124_4634_n28), .CIN(n71), .COUT(DP_OP_357J3_124_4634_n9), 
        .SUM(N386) );
  FULLADD DP_OP_357J3_124_4634_U9 ( .A(DP_OP_357J3_124_4634_n25), .B(
        DP_OP_357J3_124_4634_n26), .CIN(n68), .COUT(DP_OP_357J3_124_4634_n8), 
        .SUM(N387) );
  FULLADD DP_OP_357J3_124_4634_U8 ( .A(DP_OP_357J3_124_4634_n23), .B(
        DP_OP_357J3_124_4634_n24), .CIN(n63), .COUT(DP_OP_357J3_124_4634_n7), 
        .SUM(N388) );
  FULLADD DP_OP_357J3_124_4634_U7 ( .A(DP_OP_357J3_124_4634_n21), .B(
        DP_OP_357J3_124_4634_n22), .CIN(n70), .COUT(DP_OP_357J3_124_4634_n6), 
        .SUM(N389) );
  FULLADD DP_OP_357J3_124_4634_U6 ( .A(DP_OP_357J3_124_4634_n19), .B(
        DP_OP_357J3_124_4634_n20), .CIN(n66), .COUT(DP_OP_357J3_124_4634_n5), 
        .SUM(N390) );
  FULLADD DP_OP_357J3_124_4634_U5 ( .A(DP_OP_357J3_124_4634_n18), .B(
        DP_OP_357J3_124_4634_n17), .CIN(n67), .COUT(DP_OP_357J3_124_4634_n4), 
        .SUM(N391) );
  INVX1 DP_OP_433_158_7755_U11 ( .IN(DP_OP_433_158_7755_n38), .OUT(
        DP_OP_433_158_7755_n37) );
  NAND2X1 DP_OP_433_158_7755_U53 ( .IN1(DP_OP_433_158_7755_n69), .IN2(
        DP_OP_433_158_7755_n60), .OUT(DP_OP_433_158_7755_n33) );
  NAND3X1 U3 ( .IN1(n578), .IN2(Final_Mantissa_reg[6]), .IN3(
        Final_Mantissa_reg[5]), .OUT(n859) );
  NAND3X1 U4 ( .IN1(n483), .IN2(Multi_dataout[14]), .IN3(n623), .OUT(n470) );
  NAND3X1 U5 ( .IN1(DP_OP_433_158_7755_n1), .IN2(n198), .IN3(
        DP_OP_433_158_7755_n37), .OUT(n190) );
  NAND2X1 U6 ( .IN1(n683), .IN2(n445), .OUT(n1) );
  NOR2X1 U7 ( .IN1(n446), .IN2(n1), .OUT(n2) );
  OAI21 U8 ( .IN1(n447), .IN2(n448), .IN3(n2), .OUT(n3) );
  OAI21 U9 ( .IN1(n711), .IN2(n3), .IN3(n204), .OUT(n4) );
  NOR2X1 U10 ( .IN1(n57), .IN2(n450), .OUT(n5) );
  NAND3X1 U11 ( .IN1(n451), .IN2(n4), .IN3(n5), .OUT(n491) );
  AOI22 U12 ( .IN1(Datain1[6]), .IN2(n598), .IN3(Datain2[6]), .IN4(n595), 
        .OUT(n6) );
  OAI21 U13 ( .IN1(n599), .IN2(n600), .IN3(n6), .OUT(n7) );
  AOI21 U14 ( .IN1(n113), .IN2(n597), .IN3(n596), .OUT(n8) );
  NOR2X1 U15 ( .IN1(n7), .IN2(n8), .OUT(n9) );
  INVX1 U16 ( .IN(n9), .OUT(n601) );
  INVX1 U17 ( .IN(n448), .OUT(n10) );
  AOI21 U18 ( .IN1(n266), .IN2(n267), .IN3(n10), .OUT(n393) );
  OAI21 U19 ( .IN1(Multi_dataout[5]), .IN2(n258), .IN3(n196), .OUT(n122) );
  NAND2X1 U20 ( .IN1(DP_OP_433_158_7755_n16), .IN2(n379), .OUT(n11) );
  INVX1 U21 ( .IN(n11), .OUT(n12) );
  OAI21 U22 ( .IN1(DP_OP_433_158_7755_n1), .IN2(Final_Exponent_reg[4]), .IN3(
        n12), .OUT(n325) );
  NAND3X1 U23 ( .IN1(n449), .IN2(n447), .IN3(n688), .OUT(n646) );
  INVX1 U24 ( .IN(n102), .OUT(n13) );
  MUX2X1 U25 ( .IN1(n102), .IN2(n13), .S(n309), .OUT(n14) );
  AOI22 U26 ( .IN1(n14), .IN2(n370), .IN3(n347), .IN4(n13), .OUT(n284) );
  NAND3X1 U27 ( .IN1(n384), .IN2(n454), .IN3(n356), .OUT(n15) );
  NOR2X1 U28 ( .IN1(n360), .IN2(n15), .OUT(n16) );
  INVX1 U29 ( .IN(n428), .OUT(n17) );
  NAND3X1 U30 ( .IN1(n457), .IN2(n16), .IN3(n17), .OUT(n626) );
  NOR2X1 U31 ( .IN1(n722), .IN2(n940), .OUT(n18) );
  AOI21 U32 ( .IN1(n18), .IN2(n673), .IN3(n674), .OUT(n19) );
  INVX1 U33 ( .IN(n19), .OUT(n728) );
  AOI21 U34 ( .IN1(n577), .IN2(n110), .IN3(n861), .OUT(n20) );
  AOI22 U35 ( .IN1(n598), .IN2(Datain1[5]), .IN3(n20), .IN4(n597), .OUT(n21)
         );
  NOR2X1 U36 ( .IN1(n649), .IN2(n599), .OUT(n22) );
  AOI21 U37 ( .IN1(n595), .IN2(Datain2[5]), .IN3(n22), .OUT(n23) );
  NAND2X1 U38 ( .IN1(n21), .IN2(n23), .OUT(n579) );
  AOI21 U39 ( .IN1(DP_OP_433_158_7755_n52), .IN2(Final_Exponent_reg[5]), .IN3(
        DP_OP_433_158_7755_n13), .OUT(n24) );
  INVX1 U40 ( .IN(n24), .OUT(C276_DATA3_5) );
  INVX1 U41 ( .IN(n319), .OUT(n25) );
  NAND3X1 U42 ( .IN1(n204), .IN2(Final_Exponent_reg[4]), .IN3(n25), .OUT(n321)
         );
  INVX1 U43 ( .IN(n205), .OUT(n26) );
  NOR2X1 U44 ( .IN1(n344), .IN2(n26), .OUT(n177) );
  NAND3X1 U45 ( .IN1(n215), .IN2(n214), .IN3(n213), .OUT(n893) );
  INVX1 U46 ( .IN(n680), .OUT(n27) );
  OAI21 U47 ( .IN1(n647), .IN2(n27), .IN3(n719), .OUT(n716) );
  NAND3X1 U48 ( .IN1(n104), .IN2(n99), .IN3(StateMC[1]), .OUT(n888) );
  NAND3X1 U49 ( .IN1(n705), .IN2(Multi_dataout[14]), .IN3(n482), .OUT(n548) );
  AOI21 U50 ( .IN1(DP_OP_433_158_7755_n75), .IN2(Final_Exponent_reg[0]), .IN3(
        DP_OP_433_158_7755_n68), .OUT(n28) );
  INVX1 U51 ( .IN(n28), .OUT(C276_DATA3_0) );
  AOI21 U52 ( .IN1(DP_OP_433_158_7755_n46), .IN2(Final_Exponent_reg[6]), .IN3(
        DP_OP_433_158_7755_n10), .OUT(n29) );
  INVX1 U53 ( .IN(n29), .OUT(C276_DATA3_6) );
  AOI21 U54 ( .IN1(n668), .IN2(n695), .IN3(n179), .OUT(n30) );
  INVX1 U55 ( .IN(n30), .OUT(n194) );
  NAND3X1 U56 ( .IN1(n330), .IN2(Final_Exponent_reg[5]), .IN3(
        Final_Exponent_reg[6]), .OUT(n340) );
  NAND3X1 U57 ( .IN1(n542), .IN2(Final_Mantissa_reg[4]), .IN3(
        Final_Mantissa_reg[3]), .OUT(n577) );
  INVX1 U58 ( .IN(Mode[0]), .OUT(n31) );
  NAND3X1 U59 ( .IN1(Mode[2]), .IN2(Mode[1]), .IN3(n31), .OUT(n643) );
  NOR2X1 U60 ( .IN1(n762), .IN2(n761), .OUT(n32) );
  INVX1 U61 ( .IN(n32), .OUT(n201) );
  NOR2X1 U62 ( .IN1(n114), .IN2(Final_Mantissa_reg[0]), .OUT(n33) );
  MUX2X1 U63 ( .IN1(Final_Mantissa_reg[0]), .IN2(n33), .S(G_reg), .OUT(n34) );
  AOI22 U64 ( .IN1(n744), .IN2(n34), .IN3(n598), .IN4(Datain1[0]), .OUT(n35)
         );
  NAND2X1 U65 ( .IN1(n860), .IN2(n35), .OUT(n36) );
  AOI21 U66 ( .IN1(n595), .IN2(Datain2[0]), .IN3(n36), .OUT(n485) );
  INVX1 U67 ( .IN(DP_OP_433_158_7755_n68), .OUT(n37) );
  INVX1 U68 ( .IN(DP_OP_433_158_7755_n67), .OUT(n38) );
  NOR2X1 U69 ( .IN1(DP_OP_433_158_7755_n66), .IN2(n38), .OUT(n39) );
  MUX2X1 U70 ( .IN1(n37), .IN2(DP_OP_433_158_7755_n68), .S(n39), .OUT(
        C276_DATA3_1) );
  INVX1 U71 ( .IN(DP_OP_433_158_7755_n64), .OUT(n40) );
  INVX1 U72 ( .IN(DP_OP_433_158_7755_n63), .OUT(n41) );
  NOR2X1 U73 ( .IN1(DP_OP_433_158_7755_n62), .IN2(n41), .OUT(n42) );
  MUX2X1 U74 ( .IN1(n40), .IN2(DP_OP_433_158_7755_n64), .S(n42), .OUT(
        C276_DATA3_2) );
  AOI21 U75 ( .IN1(DP_OP_433_158_7755_n42), .IN2(Final_Exponent_reg[7]), .IN3(
        DP_OP_433_158_7755_n7), .OUT(n43) );
  INVX1 U76 ( .IN(n43), .OUT(C276_DATA3_7) );
  INVX1 U77 ( .IN(DP_OP_357J3_124_4634_n4), .OUT(n44) );
  MUX2X1 U78 ( .IN1(n44), .IN2(DP_OP_357J3_124_4634_n4), .S(n62), .OUT(N392)
         );
  OAI21 U79 ( .IN1(n55), .IN2(n855), .IN3(n851), .OUT(n164) );
  INVX1 U80 ( .IN(n725), .OUT(n45) );
  AOI22 U81 ( .IN1(n719), .IN2(n708), .IN3(Debug_reg[2]), .IN4(n715), .OUT(n46) );
  AOI22 U82 ( .IN1(n719), .IN2(n709), .IN3(n46), .IN4(n720), .OUT(n47) );
  INVX1 U83 ( .IN(n122), .OUT(n48) );
  OAI21 U84 ( .IN1(n710), .IN2(n48), .IN3(n719), .OUT(n49) );
  AOI22 U85 ( .IN1(n719), .IN2(n711), .IN3(n47), .IN4(n49), .OUT(n50) );
  NAND2X1 U86 ( .IN1(Multi_dataout[14]), .IN2(n722), .OUT(n51) );
  NOR2X1 U87 ( .IN1(n51), .IN2(n712), .OUT(n52) );
  AOI21 U88 ( .IN1(n728), .IN2(Debug_reg[2]), .IN3(n52), .OUT(n53) );
  NAND2X1 U89 ( .IN1(n45), .IN2(n727), .OUT(n54) );
  OAI21 U90 ( .IN1(n50), .IN2(n54), .IN3(n53), .OUT(n144) );
  INVX4 U91 ( .IN(Exc_Ack_BAR), .OUT(n55) );
  NAND2X1 U92 ( .IN1(Datain2[11]), .IN2(n768), .OUT(n83) );
  INVX4 U93 ( .IN(n709), .OUT(n56) );
  INVX1 U94 ( .IN(Datain2[11]), .OUT(n758) );
  NAND2X1 U95 ( .IN1(Datain1[11]), .IN2(Datain2[11]), .OUT(n85) );
  NAND2X1 U96 ( .IN1(Datain1[10]), .IN2(Datain2[10]), .OUT(n82) );
  BUF4X U97 ( .IN(n452), .OUT(n57) );
  BUF4X U98 ( .IN(n565), .OUT(n58) );
  INVX1 U99 ( .IN(n565), .OUT(n59) );
  NANDX2 U100 ( .IN1(DP_OP_433_158_7755_n1), .IN2(n227), .OUT(
        DP_OP_433_158_7755_n46) );
  BUF8X U101 ( .IN(DP_OP_433_158_7755_n56), .OUT(DP_OP_433_158_7755_n1) );
  INVX1 U102 ( .IN(Datain1[9]), .OUT(n765) );
  NANDX2 U103 ( .IN1(n318), .IN2(n317), .OUT(n877) );
  NANDX2 U104 ( .IN1(n315), .IN2(n314), .OUT(n316) );
  NANDX2 U105 ( .IN1(n308), .IN2(n317), .OUT(n878) );
  NANDX2 U106 ( .IN1(n301), .IN2(n317), .OUT(n879) );
  NAND2X1 U107 ( .IN1(n609), .IN2(n567), .OUT(n573) );
  NANDX2 U108 ( .IN1(n551), .IN2(n550), .OUT(n552) );
  NAND2X1 U109 ( .IN1(n609), .IN2(n570), .OUT(n495) );
  NANDX2 U110 ( .IN1(n306), .IN2(n305), .OUT(n307) );
  NAND2X1 U111 ( .IN1(n627), .IN2(n626), .OUT(n192) );
  INVX1 U112 ( .IN(n665), .OUT(n666) );
  NANDX2 U113 ( .IN1(n427), .IN2(n426), .OUT(n433) );
  INVX1 U114 ( .IN(n269), .OUT(n270) );
  NAND2X1 U115 ( .IN1(n374), .IN2(N391), .OUT(n375) );
  INVX1 U116 ( .IN(n354), .OUT(n355) );
  BUF4X U117 ( .IN(DP_OP_357J3_124_4634_n5), .OUT(n67) );
  NAND2X1 U118 ( .IN1(n374), .IN2(N390), .OUT(n348) );
  INVX1 U119 ( .IN(n428), .OUT(n431) );
  INVX1 U120 ( .IN(n254), .OUT(n255) );
  NANDX2 U121 ( .IN1(n279), .IN2(n399), .OUT(n281) );
  BUF4X U122 ( .IN(DP_OP_357J3_124_4634_n7), .OUT(n70) );
  INVX1 U123 ( .IN(n716), .OUT(n717) );
  NANDX2 U124 ( .IN1(n418), .IN2(n417), .OUT(n419) );
  NAND2X1 U125 ( .IN1(n374), .IN2(N387), .OUT(n285) );
  BUF4X U126 ( .IN(DP_OP_357J3_124_4634_n8), .OUT(n63) );
  INVX1 U127 ( .IN(n372), .OUT(n341) );
  NAND2X1 U128 ( .IN1(n719), .IN2(n685), .OUT(n686) );
  NAND2X1 U129 ( .IN1(n655), .IN2(n714), .OUT(n656) );
  INVX1 U130 ( .IN(n640), .OUT(n166) );
  INVX1 U131 ( .IN(n934), .OUT(n130) );
  INVX1 U132 ( .IN(n932), .OUT(n132) );
  INVX1 U133 ( .IN(n930), .OUT(n134) );
  NAND2X1 U134 ( .IN1(n676), .IN2(n675), .OUT(n677) );
  NAND2X1 U135 ( .IN1(n374), .IN2(N384), .OUT(n296) );
  INVX1 U136 ( .IN(n933), .OUT(n131) );
  NANDX2 U137 ( .IN1(n246), .IN2(n647), .OUT(n356) );
  NANDX2 U138 ( .IN1(Debug_reg[1]), .IN2(n728), .OUT(n186) );
  NAND2X1 U139 ( .IN1(n205), .IN2(n479), .OUT(n480) );
  INVX1 U140 ( .IN(n928), .OUT(n136) );
  INVX1 U141 ( .IN(n931), .OUT(n133) );
  INVX4 U142 ( .IN(n384), .OUT(n386) );
  INVX1 U143 ( .IN(n929), .OUT(n135) );
  INVX1 U144 ( .IN(n926), .OUT(n138) );
  NAND2X1 U145 ( .IN1(n205), .IN2(n620), .OUT(n621) );
  INVX1 U146 ( .IN(n927), .OUT(n137) );
  INVX1 U147 ( .IN(n924), .OUT(n140) );
  INVX1 U148 ( .IN(n935), .OUT(n129) );
  INVX1 U149 ( .IN(n938), .OUT(n128) );
  INVX1 U150 ( .IN(n923), .OUT(n141) );
  INVX1 U151 ( .IN(n740), .OUT(n850) );
  INVX1 U152 ( .IN(n925), .OUT(n139) );
  NAND2X1 U153 ( .IN1(n719), .IN2(n653), .OUT(n655) );
  INVX1 U154 ( .IN(n901), .OUT(n162) );
  INVX1 U155 ( .IN(n898), .OUT(n163) );
  BUF4X U156 ( .IN(DP_OP_357J3_124_4634_n10), .OUT(n71) );
  NAND2X1 U157 ( .IN1(n825), .IN2(n824), .OUT(n826) );
  NANDX2 U158 ( .IN1(n411), .IN2(n231), .OUT(n384) );
  NANDX2 U159 ( .IN1(T_reg), .IN2(n474), .OUT(n464) );
  NANDX2 U160 ( .IN1(G_reg), .IN2(n474), .OUT(n475) );
  INVX1 U161 ( .IN(n736), .OUT(n699) );
  INVX1 U162 ( .IN(n648), .OUT(n231) );
  NANDX2 U163 ( .IN1(Final_Exponent_reg[7]), .IN2(n371), .OUT(n220) );
  INVX1 U164 ( .IN(n339), .OUT(n342) );
  INVX1 U165 ( .IN(n843), .OUT(n881) );
  BUF4X U166 ( .IN(DP_OP_357J3_124_4634_n11), .OUT(n69) );
  INVX1 U167 ( .IN(n904), .OUT(n159) );
  INVX1 U168 ( .IN(n275), .OUT(n276) );
  INVX1 U169 ( .IN(n905), .OUT(n158) );
  INVX1 U170 ( .IN(n903), .OUT(n160) );
  INVX1 U171 ( .IN(n907), .OUT(n156) );
  INVX1 U172 ( .IN(n908), .OUT(n155) );
  INVX1 U173 ( .IN(n910), .OUT(n154) );
  INVX1 U174 ( .IN(n911), .OUT(n153) );
  INVX1 U175 ( .IN(n906), .OUT(n157) );
  INVX1 U176 ( .IN(n902), .OUT(n161) );
  NAND2X1 U177 ( .IN1(n146), .IN2(n894), .OUT(n143) );
  INVX1 U178 ( .IN(n918), .OUT(n147) );
  INVX1 U179 ( .IN(n916), .OUT(n148) );
  INVX1 U180 ( .IN(n915), .OUT(n149) );
  INVX1 U181 ( .IN(n913), .OUT(n151) );
  INVX1 U182 ( .IN(n914), .OUT(n150) );
  INVX1 U183 ( .IN(n912), .OUT(n152) );
  INVX4 U184 ( .IN(Multi_ack), .OUT(n750) );
  NAND2X1 U185 ( .IN1(n623), .IN2(Multi_dataout[15]), .OUT(n459) );
  NANDX2 U186 ( .IN1(n413), .IN2(n256), .OUT(n421) );
  INVX1 U187 ( .IN(n783), .OUT(n788) );
  NAND2X1 U188 ( .IN1(n747), .IN2(n853), .OUT(n637) );
  NAND2X1 U189 ( .IN1(n747), .IN2(n854), .OUT(n633) );
  NAND2X1 U190 ( .IN1(n482), .IN2(Multi_dataout[15]), .OUT(n275) );
  INVX1 U191 ( .IN(n789), .OUT(Dataout[15]) );
  INVX1 U192 ( .IN(n817), .OUT(Exc[2]) );
  NANDX2 U193 ( .IN1(n98), .IN2(n398), .OUT(n246) );
  NANDX2 U194 ( .IN1(n319), .IN2(n262), .OUT(n261) );
  NAND2X1 U195 ( .IN1(n940), .IN2(n939), .OUT(n849) );
  INVX1 U196 ( .IN(n895), .OUT(n351) );
  NANDX2 U197 ( .IN1(n413), .IN2(n260), .OUT(n262) );
  NANDX2 U198 ( .IN1(n108), .IN2(Dataout_valid), .OUT(n817) );
  NANDX2 U199 ( .IN1(Final_Mantissa_reg[2]), .IN2(n222), .OUT(n541) );
  NAND2X1 U200 ( .IN1(n55), .IN2(n852), .OUT(n778) );
  NAND2X1 U201 ( .IN1(n812), .IN2(n55), .OUT(n634) );
  NAND2X1 U202 ( .IN1(n845), .IN2(n205), .OUT(n848) );
  INVX1 U203 ( .IN(n858), .OUT(n277) );
  INVX1 U204 ( .IN(n793), .OUT(Debug[4]) );
  INVX1 U205 ( .IN(n730), .OUT(Debug[3]) );
  INVX1 U206 ( .IN(n713), .OUT(Debug[2]) );
  INVX1 U207 ( .IN(n672), .OUT(Debug[0]) );
  INVX1 U208 ( .IN(n704), .OUT(Debug[1]) );
  NANDX2 U209 ( .IN1(Final_Exponent_reg[3]), .IN2(n310), .OUT(n319) );
  NANDX2 U210 ( .IN1(n98), .IN2(n266), .OUT(n260) );
  NAND2X1 U211 ( .IN1(n891), .IN2(n810), .OUT(n812) );
  INVX1 U212 ( .IN(n854), .OUT(n852) );
  INVX1 U213 ( .IN(n631), .OUT(n890) );
  NANDX2 U214 ( .IN1(Datain1[12]), .IN2(n88), .OUT(n87) );
  NANDX2 U215 ( .IN1(Final_Mantissa_reg[1]), .IN2(n221), .OUT(n522) );
  NANDX2 U216 ( .IN1(Datain1[11]), .IN2(n758), .OUT(n84) );
  NANDX2 U217 ( .IN1(Datain1[13]), .IN2(n93), .OUT(n91) );
  NANDX2 U218 ( .IN1(StateMC[0]), .IN2(n743), .OUT(n821) );
  NANDX2 U219 ( .IN1(StateMC[0]), .IN2(n223), .OUT(n820) );
  NAND2X1 U220 ( .IN1(n205), .IN2(n884), .OUT(n939) );
  INVX1 U221 ( .IN(DP_OP_357J3_124_4634_n15), .OUT(n62) );
  NANDX2 U222 ( .IN1(Datain1[13]), .IN2(Datain2[13]), .OUT(n95) );
  NANDX2 U223 ( .IN1(Datain1[12]), .IN2(Datain2[12]), .OUT(n89) );
  INVX1 U224 ( .IN(n504), .OUT(n221) );
  NANDX2 U225 ( .IN1(DP_OP_357J3_124_4634_n66), .IN2(DP_OP_357J3_124_4634_n58), 
        .OUT(n74) );
  NANDX2 U226 ( .IN1(n101), .IN2(n114), .OUT(n632) );
  NANDX2 U227 ( .IN1(StateMC[2]), .IN2(StateMC[1]), .OUT(n224) );
  INVX4 U228 ( .IN(DP_OP_357J3_124_4634_n66), .OUT(n60) );
  INVX4 U229 ( .IN(DP_OP_357J3_124_4634_n58), .OUT(n61) );
  NANDX2 U230 ( .IN1(n99), .IN2(n105), .OUT(n884) );
  NANDX2 U231 ( .IN1(Mode[2]), .IN2(Mode[0]), .OUT(n732) );
  NANDX2 U232 ( .IN1(n104), .IN2(n743), .OUT(n810) );
  INVX1 U233 ( .IN(Datain2[13]), .OUT(n93) );
  INVX1 U234 ( .IN(Datain1[13]), .OUT(n92) );
  NAND2X1 U235 ( .IN1(Datain2[13]), .IN2(n92), .OUT(n90) );
  INVX1 U236 ( .IN(Datain2[12]), .OUT(n88) );
  NAND2X1 U237 ( .IN1(Datain2[12]), .IN2(n767), .OUT(n86) );
  INVX1 U238 ( .IN(Datain1[10]), .OUT(n81) );
  NAND2X1 U239 ( .IN1(Datain2[10]), .IN2(n81), .OUT(n79) );
  INVX1 U240 ( .IN(Datain2[9]), .OUT(n77) );
  NAND2X1 U241 ( .IN1(DP_OP_357J3_124_4634_n66), .IN2(n61), .OUT(n73) );
  NAND2X1 U242 ( .IN1(DP_OP_357J3_124_4634_n58), .IN2(n60), .OUT(n72) );
  INVX4 U243 ( .IN(n95), .OUT(DP_OP_357J3_124_4634_n18) );
  NANDX2 U244 ( .IN1(n91), .IN2(n90), .OUT(DP_OP_357J3_124_4634_n19) );
  INVX4 U245 ( .IN(n89), .OUT(DP_OP_357J3_124_4634_n20) );
  NANDX2 U246 ( .IN1(n87), .IN2(n86), .OUT(DP_OP_357J3_124_4634_n21) );
  INVX4 U247 ( .IN(n85), .OUT(DP_OP_357J3_124_4634_n22) );
  NANDX2 U248 ( .IN1(n84), .IN2(n83), .OUT(DP_OP_357J3_124_4634_n23) );
  INVX4 U249 ( .IN(n82), .OUT(DP_OP_357J3_124_4634_n24) );
  NANDX2 U250 ( .IN1(n80), .IN2(n79), .OUT(DP_OP_357J3_124_4634_n25) );
  INVX4 U251 ( .IN(n78), .OUT(DP_OP_357J3_124_4634_n26) );
  NANDX2 U252 ( .IN1(n76), .IN2(n75), .OUT(DP_OP_357J3_124_4634_n27) );
  INVX4 U253 ( .IN(n74), .OUT(DP_OP_357J3_124_4634_n28) );
  INVX4 U254 ( .IN(RSOP_428_C1_Z_0), .OUT(n65) );
  NANDX2 U255 ( .IN1(n73), .IN2(n72), .OUT(DP_OP_357J3_124_4634_n29) );
  NAND2X1 U256 ( .IN1(Datain1[10]), .IN2(n757), .OUT(n80) );
  NAND2X1 U257 ( .IN1(Datain2[9]), .IN2(n765), .OUT(n75) );
  NAND2X1 U258 ( .IN1(Datain1[9]), .IN2(Datain2[9]), .OUT(n78) );
  NAND2X1 U259 ( .IN1(Datain1[9]), .IN2(n77), .OUT(n76) );
  BUF4X U260 ( .IN(DP_OP_357J3_124_4634_n6), .OUT(n66) );
  BUF4X U261 ( .IN(DP_OP_357J3_124_4634_n9), .OUT(n68) );
  NAND2X1 U262 ( .IN1(n379), .IN2(C276_DATA3_2), .OUT(n314) );
  INVX1 U263 ( .IN(n127), .OUT(N90) );
  NAND2X1 U264 ( .IN1(n416), .IN2(n647), .OUT(n404) );
  NANDX2 U265 ( .IN1(n810), .IN2(n861), .OUT(n212) );
  NANDX2 U266 ( .IN1(n191), .IN2(n190), .OUT(n628) );
  NAND2X1 U267 ( .IN1(n197), .IN2(DP_OP_433_158_7755_n56), .OUT(n198) );
  NANDX2 U268 ( .IN1(n740), .IN2(n741), .OUT(n183) );
  NANDX2 U269 ( .IN1(n727), .IN2(Multi_ack), .OUT(n712) );
  NANDX2 U270 ( .IN1(n850), .IN2(n481), .OUT(n599) );
  INVX4 U271 ( .IN(Multi_dataout[10]), .OUT(n586) );
  INVX4 U272 ( .IN(n857), .OUT(n477) );
  NANDX2 U273 ( .IN1(n586), .IN2(n232), .OUT(n233) );
  NANDX2 U274 ( .IN1(n390), .IN2(n451), .OUT(n392) );
  INVX4 U275 ( .IN(n643), .OUT(n644) );
  NANDX2 U276 ( .IN1(n204), .IN2(n310), .OUT(n309) );
  NAND2X1 U277 ( .IN1(Final_Exponent_reg[0]), .IN2(Final_Exponent_reg[1]), 
        .OUT(n244) );
  NANDX2 U278 ( .IN1(Multi_dataout[0]), .IN2(n603), .OUT(n466) );
  NAND2X1 U279 ( .IN1(n623), .IN2(n622), .OUT(n624) );
  NANDX2 U280 ( .IN1(n363), .IN2(n430), .OUT(C1_Z_1) );
  NAND2X1 U281 ( .IN1(n122), .IN2(n692), .OUT(n659) );
  NANDX2 U282 ( .IN1(n744), .IN2(n859), .OUT(n596) );
  NANDX2 U283 ( .IN1(n732), .IN2(n643), .OUT(n792) );
  NANDX2 U284 ( .IN1(n939), .IN2(n642), .OUT(n474) );
  NANDX2 U285 ( .IN1(n483), .IN2(n742), .OUT(n484) );
  NANDX2 U286 ( .IN1(n205), .IN2(n194), .OUT(n193) );
  NANDX2 U287 ( .IN1(n421), .IN2(n420), .OUT(n445) );
  NAND2X1 U288 ( .IN1(n719), .IN2(n658), .OUT(n720) );
  NANDX2 U289 ( .IN1(n644), .IN2(n746), .OUT(n737) );
  NANDX2 U290 ( .IN1(n178), .IN2(N392), .OUT(n175) );
  INVX4 U291 ( .IN(n452), .OUT(n357) );
  NANDX2 U292 ( .IN1(n413), .IN2(n397), .OUT(n454) );
  INVX4 U293 ( .IN(Multi_dataout[15]), .OUT(n483) );
  NAND2X1 U294 ( .IN1(Final_Mantissa_reg[0]), .IN2(G_reg), .OUT(n504) );
  BUF4X U295 ( .IN(n937), .OUT(n203) );
  NANDX2 U296 ( .IN1(n167), .IN2(n165), .OUT(n883) );
  NANDX2 U297 ( .IN1(n195), .IN2(n193), .OUT(n94) );
  NANDX2 U298 ( .IN1(n183), .IN2(n180), .OUT(n179) );
  INVX4 U299 ( .IN(n889), .OUT(n745) );
  NANDX2 U300 ( .IN1(n483), .IN2(n282), .OUT(n622) );
  NANDX2 U301 ( .IN1(n471), .IN2(n250), .OUT(n237) );
  NANDX2 U302 ( .IN1(n808), .IN2(n55), .OUT(n851) );
  BUF4X U303 ( .IN(n917), .OUT(n202) );
  NANDX2 U304 ( .IN1(n205), .IN2(n738), .OUT(n739) );
  NANDX2 U305 ( .IN1(n185), .IN2(n200), .OUT(n184) );
  INVX1 U306 ( .IN(n688), .OUT(n709) );
  INVX4 U307 ( .IN(n237), .OUT(n174) );
  INVX4 U308 ( .IN(Multi_dataout[8]), .OUT(n537) );
  INVX4 U309 ( .IN(n851), .OUT(n273) );
  NANDX2 U310 ( .IN1(n205), .IN2(n292), .OUT(n200) );
  INVX4 U311 ( .IN(n840), .OUT(n909) );
  INVX4 U312 ( .IN(Datain1[12]), .OUT(n767) );
  INVX1 U313 ( .IN(n201), .OUT(n841) );
  INVX4 U314 ( .IN(Datain2[10]), .OUT(n757) );
  INVX1 U315 ( .IN(n810), .OUT(n784) );
  INVX4 U316 ( .IN(n739), .OUT(n96) );
  NANDX2 U317 ( .IN1(n611), .IN2(n567), .OUT(n496) );
  NAND2X1 U318 ( .IN1(n692), .IN2(n449), .OUT(n711) );
  NANDX2 U319 ( .IN1(n442), .IN2(n439), .OUT(n437) );
  NANDX2 U320 ( .IN1(n439), .IN2(n438), .OUT(n440) );
  INVX4 U321 ( .IN(n212), .OUT(n217) );
  NAND2X1 U322 ( .IN1(n652), .IN2(n651), .OUT(n653) );
  NANDX2 U323 ( .IN1(n448), .IN2(n265), .OUT(n271) );
  INVX4 U324 ( .IN(n421), .OUT(n259) );
  NAND2X1 U325 ( .IN1(n243), .IN2(n684), .OUT(n651) );
  INVX4 U326 ( .IN(n401), .OUT(n241) );
  INVX4 U327 ( .IN(n659), .OUT(n280) );
  INVX4 U328 ( .IN(n126), .OUT(n123) );
  NANDX2 U329 ( .IN1(n196), .IN2(n688), .OUT(n126) );
  NANDX2 U330 ( .IN1(n683), .IN2(n174), .OUT(n173) );
  NANDX2 U331 ( .IN1(n569), .IN2(n537), .OUT(n234) );
  NANDX2 U332 ( .IN1(n649), .IN2(n565), .OUT(n230) );
  NANDX2 U333 ( .IN1(n291), .IN2(n290), .OUT(n370) );
  NANDX2 U334 ( .IN1(n273), .IN2(n854), .OUT(n561) );
  NANDX2 U335 ( .IN1(n181), .IN2(n180), .OUT(n292) );
  NANDX2 U336 ( .IN1(n201), .IN2(n909), .OUT(n207) );
  INVX4 U337 ( .IN(Datain2[7]), .OUT(n760) );
  INVX4 U338 ( .IN(n897), .OUT(n899) );
  NANDX2 U339 ( .IN1(n205), .IN2(n750), .OUT(n920) );
  NANDX2 U340 ( .IN1(n706), .IN2(n705), .OUT(n725) );
  NANDX2 U341 ( .IN1(n533), .IN2(n532), .OUT(n534) );
  NANDX2 U342 ( .IN1(n609), .IN2(n518), .OUT(n533) );
  NANDX2 U343 ( .IN1(n515), .IN2(n514), .OUT(n516) );
  NANDX2 U344 ( .IN1(n609), .IN2(n587), .OUT(n515) );
  NANDX2 U345 ( .IN1(n545), .IN2(n544), .OUT(n546) );
  INVX4 U346 ( .IN(n599), .OUT(n547) );
  NANDX2 U347 ( .IN1(n494), .IN2(n493), .OUT(n570) );
  NANDX2 U348 ( .IN1(n490), .IN2(n489), .OUT(n567) );
  INVX4 U349 ( .IN(n636), .OUT(n835) );
  NANDX2 U350 ( .IN1(n501), .IN2(n500), .OUT(n587) );
  INVX4 U351 ( .IN(n538), .OUT(n588) );
  NANDX2 U352 ( .IN1(n613), .IN2(n611), .OUT(n538) );
  NANDX2 U353 ( .IN1(n503), .IN2(n502), .OUT(n582) );
  NANDX2 U354 ( .IN1(n520), .IN2(n519), .OUT(n608) );
  NANDX2 U355 ( .IN1(n675), .IN2(n491), .OUT(n492) );
  NANDX2 U356 ( .IN1(n607), .IN2(n606), .OUT(n610) );
  INVX4 U357 ( .IN(n549), .OUT(n611) );
  INVX4 U358 ( .IN(n484), .OUT(n705) );
  NANDX2 U359 ( .IN1(n675), .IN2(n488), .OUT(n549) );
  NANDX2 U360 ( .IN1(n895), .IN2(n480), .OUT(n618) );
  NANDX2 U361 ( .IN1(n700), .IN2(n701), .OUT(n189) );
  NANDX2 U362 ( .IN1(n694), .IN2(n693), .OUT(n700) );
  NANDX2 U363 ( .IN1(n722), .IN2(n695), .OUT(n736) );
  NANDX2 U364 ( .IN1(n458), .IN2(n457), .OUT(n613) );
  NANDX2 U365 ( .IN1(n444), .IN2(n443), .OUT(n518) );
  INVX4 U366 ( .IN(n491), .OUT(n488) );
  NANDX2 U367 ( .IN1(n468), .IN2(n467), .OUT(n553) );
  INVX4 U368 ( .IN(n437), .OUT(n605) );
  NANDX2 U369 ( .IN1(n466), .IN2(n465), .OUT(n539) );
  INVX4 U370 ( .IN(n581), .OUT(n521) );
  NANDX2 U371 ( .IN1(n438), .IN2(n441), .OUT(n581) );
  INVX4 U372 ( .IN(n440), .OUT(n604) );
  INVX4 U373 ( .IN(n442), .OUT(n438) );
  INVX4 U374 ( .IN(n441), .OUT(n439) );
  INVX4 U375 ( .IN(n585), .OUT(n603) );
  NANDX2 U376 ( .IN1(n442), .IN2(n441), .OUT(n585) );
  NANDX2 U377 ( .IN1(n410), .IN2(n409), .OUT(n442) );
  NANDX2 U378 ( .IN1(n422), .IN2(n402), .OUT(n446) );
  NANDX2 U379 ( .IN1(n398), .IN2(n397), .OUT(n422) );
  INVX4 U380 ( .IN(n389), .OUT(n451) );
  NANDX2 U381 ( .IN1(n388), .IN2(n387), .OUT(n389) );
  NANDX2 U382 ( .IN1(n217), .IN2(n216), .OUT(n781) );
  NANDX2 U383 ( .IN1(n634), .IN2(n633), .OUT(n636) );
  INVX4 U384 ( .IN(n224), .OUT(n743) );
  INVX4 U385 ( .IN(n632), .OUT(n823) );
  NANDX2 U386 ( .IN1(n629), .IN2(n628), .OUT(n668) );
  INVX4 U387 ( .IN(n459), .OUT(n625) );
  NANDX2 U388 ( .IN1(n645), .IN2(n719), .OUT(n676) );
  NANDX2 U389 ( .IN1(n642), .IN2(n641), .OUT(n674) );
  NANDX2 U390 ( .IN1(n727), .IN2(n750), .OUT(n642) );
  NANDX2 U391 ( .IN1(n176), .IN2(n175), .OUT(n380) );
  INVX4 U392 ( .IN(n370), .OUT(n332) );
  INVX4 U393 ( .IN(n184), .OUT(n352) );
  NANDX2 U394 ( .IN1(n200), .IN2(n329), .OUT(n875) );
  NANDX2 U395 ( .IN1(n359), .IN2(n387), .OUT(n368) );
  NANDX2 U396 ( .IN1(n366), .IN2(n356), .OUT(n450) );
  INVX4 U397 ( .IN(C1_Z_3), .OUT(n199) );
  NANDX2 U398 ( .IN1(n675), .IN2(n626), .OUT(n272) );
  NANDX2 U399 ( .IN1(n271), .IN2(n429), .OUT(n452) );
  NANDX2 U400 ( .IN1(n393), .IN2(n678), .OUT(n429) );
  INVX4 U401 ( .IN(n449), .OUT(n678) );
  INVX4 U402 ( .IN(n262), .OUT(n448) );
  NANDX2 U403 ( .IN1(n361), .IN2(n430), .OUT(n391) );
  NANDX2 U404 ( .IN1(n261), .IN2(n710), .OUT(n430) );
  INVX4 U405 ( .IN(n447), .OUT(n710) );
  NANDX2 U406 ( .IN1(n259), .IN2(n420), .OUT(n361) );
  INVX4 U407 ( .IN(n679), .OUT(n420) );
  NANDX2 U408 ( .IN1(n455), .IN2(n255), .OUT(n428) );
  NANDX2 U409 ( .IN1(n252), .IN2(n658), .OUT(n387) );
  NANDX2 U410 ( .IN1(n309), .IN2(n398), .OUT(n252) );
  NANDX2 U411 ( .IN1(n249), .IN2(n654), .OUT(n366) );
  INVX4 U412 ( .IN(n395), .OUT(n249) );
  NANDX2 U413 ( .IN1(n247), .IN2(n246), .OUT(n395) );
  NANDX2 U414 ( .IN1(n267), .IN2(n398), .OUT(n247) );
  INVX4 U415 ( .IN(n245), .OUT(n267) );
  NANDX2 U416 ( .IN1(n241), .IN2(n709), .OUT(n455) );
  INVX4 U417 ( .IN(n687), .OUT(n397) );
  INVX4 U418 ( .IN(n246), .OUT(n416) );
  INVX4 U419 ( .IN(n413), .OUT(n398) );
  NANDX2 U420 ( .IN1(n102), .IN2(n266), .OUT(n413) );
  INVX4 U421 ( .IN(n229), .OUT(n266) );
  INVX4 U422 ( .IN(n731), .OUT(n675) );
  NANDX2 U423 ( .IN1(n695), .IN2(n627), .OUT(n731) );
  INVX4 U424 ( .IN(n673), .OUT(n627) );
  NANDX2 U425 ( .IN1(n483), .IN2(n226), .OUT(n673) );
  INVX4 U426 ( .IN(n894), .OUT(n695) );
  NANDX2 U427 ( .IN1(n482), .IN2(Multi_ack), .OUT(n894) );
  NANDX2 U428 ( .IN1(n280), .IN2(n426), .OUT(n734) );
  INVX4 U429 ( .IN(n646), .OUT(n426) );
  NANDX2 U430 ( .IN1(n692), .IN2(n270), .OUT(n449) );
  NANDX2 U431 ( .IN1(n264), .IN2(n447), .OUT(n692) );
  NANDX2 U432 ( .IN1(Multi_dataout[2]), .IN2(n268), .OUT(n447) );
  INVX4 U433 ( .IN(n263), .OUT(n268) );
  NANDX2 U434 ( .IN1(n123), .IN2(n122), .OUT(n263) );
  NANDX2 U435 ( .IN1(n172), .IN2(n169), .OUT(n688) );
  INVX4 U436 ( .IN(n170), .OUT(n169) );
  NANDX2 U437 ( .IN1(n240), .IN2(n680), .OUT(n170) );
  INVX4 U438 ( .IN(n171), .OUT(n196) );
  NANDX2 U439 ( .IN1(n680), .IN2(n172), .OUT(n171) );
  INVX4 U440 ( .IN(n173), .OUT(n172) );
  NANDX2 U441 ( .IN1(n235), .IN2(n683), .OUT(n680) );
  NANDX2 U442 ( .IN1(n234), .IN2(n250), .OUT(n683) );
  INVX4 U443 ( .IN(n707), .OUT(n250) );
  NANDX2 U444 ( .IN1(n684), .IN2(n681), .OUT(n707) );
  INVX4 U445 ( .IN(Multi_dataout[9]), .OUT(n569) );
  NANDX2 U446 ( .IN1(n684), .IN2(n233), .OUT(n681) );
  INVX4 U447 ( .IN(n230), .OUT(n684) );
  INVX4 U448 ( .IN(Multi_dataout[13]), .OUT(n649) );
  INVX4 U449 ( .IN(n290), .OUT(n481) );
  NANDX2 U450 ( .IN1(n742), .IN2(n276), .OUT(n290) );
  INVX4 U451 ( .IN(n476), .OUT(n742) );
  NANDX2 U452 ( .IN1(n623), .IN2(Multi_ack), .OUT(n476) );
  INVX4 U453 ( .IN(n893), .OUT(n623) );
  NANDX2 U454 ( .IN1(n633), .IN2(n637), .OUT(n595) );
  INVX4 U455 ( .IN(n561), .OUT(n598) );
  INVX4 U456 ( .IN(n891), .OUT(n808) );
  NANDX2 U457 ( .IN1(n205), .IN2(n225), .OUT(n895) );
  NAND2X1 U458 ( .IN1(n104), .IN2(n223), .OUT(n631) );
  INVX4 U459 ( .IN(n884), .OUT(n223) );
  NANDX2 U460 ( .IN1(n374), .IN2(N392), .OUT(n180) );
  INVX4 U461 ( .IN(n207), .OUT(RSOP_428_C1_Z_0) );
  NANDX2 U462 ( .IN1(n746), .IN2(n218), .OUT(n825) );
  INVX4 U463 ( .IN(n833), .OUT(n218) );
  INVX4 U464 ( .IN(Datain1[11]), .OUT(n768) );
  INVX4 U465 ( .IN(n182), .OUT(n181) );
  NANDX2 U466 ( .IN1(n860), .IN2(n183), .OUT(n182) );
  INVX4 U467 ( .IN(n291), .OUT(n741) );
  NANDX2 U468 ( .IN1(n744), .IN2(n274), .OUT(n291) );
  INVX4 U469 ( .IN(n859), .OUT(n274) );
  INVX4 U470 ( .IN(n577), .OUT(n578) );
  INVX4 U471 ( .IN(n541), .OUT(n542) );
  INVX4 U472 ( .IN(n522), .OUT(n222) );
  INVX4 U473 ( .IN(n861), .OUT(n744) );
  NAND2X1 U474 ( .IN1(StateMC[0]), .IN2(n211), .OUT(n861) );
  INVX4 U475 ( .IN(n340), .OUT(n371) );
  INVX4 U476 ( .IN(n321), .OUT(n330) );
  INVX4 U477 ( .IN(n244), .OUT(n310) );
  NANDX2 U478 ( .IN1(n816), .IN2(n747), .OUT(n860) );
  NANDX2 U479 ( .IN1(n55), .IN2(n748), .OUT(n219) );
  NAND2X1 U480 ( .IN1(n104), .IN2(n211), .OUT(n855) );
  INVX4 U481 ( .IN(n206), .OUT(n211) );
  NAND2X1 U482 ( .IN1(StateMC[2]), .IN2(n105), .OUT(n206) );
  INVX4 U483 ( .IN(RSTn_BAR), .OUT(n205) );
  NAND2X1 U484 ( .IN1(Final_Exponent_reg[8]), .IN2(n630), .OUT(n195) );
  NAND2X1 U485 ( .IN1(Debug_reg[3]), .IN2(n792), .OUT(n730) );
  INVX1 U486 ( .IN(Mode[0]), .OUT(n749) );
  INVX1 U487 ( .IN(n729), .OUT(n145) );
  NAND2X1 U488 ( .IN1(n379), .IN2(C276_DATA3_1), .OUT(n305) );
  INVX1 U489 ( .IN(n299), .OUT(n300) );
  NAND2X1 U490 ( .IN1(n103), .IN2(n370), .OUT(n295) );
  INVX1 U491 ( .IN(n535), .OUT(n869) );
  NAND2X1 U492 ( .IN1(n109), .IN2(n522), .OUT(n523) );
  INVX1 U493 ( .IN(Datain1[2]), .OUT(n525) );
  INVX1 U494 ( .IN(n499), .OUT(n871) );
  INVX1 U495 ( .IN(n517), .OUT(n870) );
  NAND2X1 U496 ( .IN1(n111), .IN2(n504), .OUT(n505) );
  INVX1 U497 ( .IN(Datain1[1]), .OUT(n507) );
  NAND2X1 U498 ( .IN1(Multi_dataout[0]), .IN2(n521), .OUT(n512) );
  INVX1 U499 ( .IN(n557), .OUT(n868) );
  NAND2X1 U500 ( .IN1(n555), .IN2(n554), .OUT(n556) );
  NAND2X1 U501 ( .IN1(Multi_dataout[10]), .IN2(n602), .OUT(n550) );
  NAND2X1 U502 ( .IN1(Datain2[3]), .IN2(n595), .OUT(n544) );
  INVX1 U503 ( .IN(n576), .OUT(n867) );
  NAND2X1 U504 ( .IN1(n112), .IN2(n558), .OUT(n559) );
  NAND2X1 U505 ( .IN1(Final_Mantissa_reg[3]), .IN2(n542), .OUT(n558) );
  INVX1 U506 ( .IN(Datain1[4]), .OUT(n562) );
  INVX1 U507 ( .IN(n210), .OUT(n882) );
  INVX1 U508 ( .IN(Exc_value[1]), .OUT(n638) );
  INVX1 U509 ( .IN(n594), .OUT(n866) );
  NAND2X1 U510 ( .IN1(Multi_dataout[0]), .IN2(n613), .OUT(n580) );
  INVX1 U511 ( .IN(n619), .OUT(n865) );
  NAND2X1 U512 ( .IN1(Final_Mantissa_reg[5]), .IN2(n578), .OUT(n597) );
  NAND2X1 U513 ( .IN1(Debug_reg[1]), .IN2(n686), .OUT(n690) );
  NAND2X1 U514 ( .IN1(n697), .IN2(n696), .OUT(n698) );
  NAND2X1 U515 ( .IN1(n455), .IN2(n454), .OUT(n456) );
  INVX1 U516 ( .IN(Multi_dataout[0]), .OUT(n434) );
  INVX1 U517 ( .IN(n424), .OUT(n405) );
  INVX4 U518 ( .IN(n821), .OUT(Dataout_valid) );
  INVX1 U519 ( .IN(n811), .OUT(n814) );
  INVX1 U520 ( .IN(n671), .OUT(n863) );
  NAND2X1 U521 ( .IN1(n719), .IN2(n654), .OUT(n714) );
  NAND2X1 U522 ( .IN1(n719), .IN2(n646), .OUT(n663) );
  INVX4 U523 ( .IN(n732), .OUT(n719) );
  INVX1 U524 ( .IN(Mode[1]), .OUT(n645) );
  NAND2X1 U525 ( .IN1(n293), .IN2(n317), .OUT(n876) );
  INVX1 U526 ( .IN(n288), .OUT(n289) );
  NAND2X1 U527 ( .IN1(n371), .IN2(n370), .OUT(n373) );
  INVX1 U528 ( .IN(n335), .OUT(n336) );
  NAND2X1 U529 ( .IN1(Final_Exponent_reg[6]), .IN2(n351), .OUT(n185) );
  NAND2X1 U530 ( .IN1(n349), .IN2(n348), .OUT(n350) );
  NAND2X1 U531 ( .IN1(n340), .IN2(n370), .OUT(n372) );
  NAND2X1 U532 ( .IN1(Final_Exponent_reg[5]), .IN2(n330), .OUT(n339) );
  INVX1 U533 ( .IN(n360), .OUT(n388) );
  INVX1 U534 ( .IN(n364), .OUT(n365) );
  INVX1 U535 ( .IN(n385), .OUT(n359) );
  NAND2X1 U536 ( .IN1(n258), .IN2(n196), .OUT(n679) );
  NAND2X1 U537 ( .IN1(Multi_dataout[8]), .IN2(n569), .OUT(n248) );
  NAND2X1 U538 ( .IN1(n97), .IN2(n103), .OUT(n245) );
  INVX1 U539 ( .IN(n411), .OUT(n242) );
  NAND2X1 U540 ( .IN1(n97), .IN2(n238), .OUT(n256) );
  INVX1 U541 ( .IN(n260), .OUT(n238) );
  NAND2X1 U542 ( .IN1(Multi_dataout[5]), .IN2(n196), .OUT(n687) );
  NAND2X1 U543 ( .IN1(n97), .IN2(n416), .OUT(n411) );
  NAND2X1 U544 ( .IN1(Final_Exponent_reg[4]), .IN2(n347), .OUT(n326) );
  INVX1 U545 ( .IN(n294), .OUT(n347) );
  INVX1 U546 ( .IN(Multi_dataout[14]), .OUT(n600) );
  INVX1 U547 ( .IN(Multi_dataout[4]), .OUT(n239) );
  INVX1 U548 ( .IN(Multi_dataout[1]), .OUT(n435) );
  INVX1 U549 ( .IN(Multi_dataout[6]), .OUT(n471) );
  NAND2X1 U550 ( .IN1(Multi_dataout[3]), .IN2(n461), .OUT(n257) );
  INVX1 U551 ( .IN(Multi_dataout[5]), .OUT(n461) );
  INVX1 U552 ( .IN(n658), .OUT(n399) );
  NAND2X1 U553 ( .IN1(Multi_dataout[6]), .IN2(n250), .OUT(n251) );
  NAND2X1 U554 ( .IN1(n683), .IN2(n680), .OUT(n708) );
  INVX1 U555 ( .IN(Multi_dataout[7]), .OUT(n486) );
  NAND2X1 U556 ( .IN1(n740), .IN2(n481), .OUT(n344) );
  NAND2X1 U557 ( .IN1(n224), .IN2(n631), .OUT(n225) );
  INVX4 U558 ( .IN(n855), .OUT(n748) );
  BUF4X U559 ( .IN(Final_Exponent_reg[2]), .OUT(n204) );
  OAI21 U560 ( .IN1(n143), .IN2(n781), .IN3(n205), .OUT(n127) );
  AOI21 U561 ( .IN1(n856), .IN2(n748), .IN3(n164), .OUT(n146) );
  OAI21 U562 ( .IN1(n166), .IN2(n179), .IN3(n205), .OUT(n165) );
  AOI21 U563 ( .IN1(n120), .IN2(n830), .IN3(n168), .OUT(n167) );
  NOR2X1 U564 ( .IN1(n940), .IN2(n831), .OUT(n168) );
  AOI21 U565 ( .IN1(n178), .IN2(n182), .IN3(n177), .OUT(n176) );
  AOI21 U566 ( .IN1(n181), .IN2(n825), .IN3(RSTn_BAR), .OUT(n178) );
  OAI21 U567 ( .IN1(RSTn_BAR), .IN2(n187), .IN3(n186), .OUT(n862) );
  AOI21 U568 ( .IN1(n698), .IN2(n699), .IN3(n188), .OUT(n187) );
  OAI21 U569 ( .IN1(n737), .IN2(n702), .IN3(n189), .OUT(n188) );
  AOI21 U570 ( .IN1(n198), .IN2(n119), .IN3(n192), .OUT(n191) );
  TIEHI U571 ( .OUT(n64) );
  NOR2X1 U572 ( .IN1(Final_Exponent_reg[8]), .IN2(DP_OP_433_158_7755_n38), 
        .OUT(n197) );
  NAND2X1 U573 ( .IN1(n649), .IN2(n648), .OUT(n650) );
  NAND2X1 U574 ( .IN1(n396), .IN2(n679), .OUT(n403) );
  NAND2X1 U575 ( .IN1(n684), .IN2(n683), .OUT(n685) );
  NAND2X1 U576 ( .IN1(n719), .IN2(n707), .OUT(n715) );
  NAND2X1 U577 ( .IN1(n652), .IN2(n681), .OUT(n278) );
  INVX1 U578 ( .IN(n681), .OUT(n394) );
  BUF4X U579 ( .IN(Datain2[8]), .OUT(DP_OP_357J3_124_4634_n58) );
  BUF4X U580 ( .IN(Datain1[7]), .OUT(DP_OP_357J3_124_4634_n65) );
  NAND2X1 U581 ( .IN1(n56), .IN2(n687), .OUT(n689) );
  NAND2X1 U582 ( .IN1(n680), .IN2(n399), .OUT(n400) );
  INVX1 U583 ( .IN(n680), .OUT(n414) );
  BUF4X U584 ( .IN(Datain1[8]), .OUT(DP_OP_357J3_124_4634_n66) );
  INVX1 U585 ( .IN(n692), .OUT(n265) );
  NAND2X1 U586 ( .IN1(Multi_dataout[12]), .IN2(n649), .OUT(n652) );
  INVX1 U587 ( .IN(Multi_dataout[12]), .OUT(n565) );
  INVX1 U588 ( .IN(N392), .OUT(n702) );
  NAND2X1 U589 ( .IN1(Multi_dataout[11]), .IN2(n603), .OUT(n607) );
  INVX1 U590 ( .IN(DP_OP_433_158_7755_n59), .OUT(DP_OP_433_158_7755_n69) );
  NAND2X1 U591 ( .IN1(n684), .IN2(Multi_dataout[11]), .OUT(n648) );
  INVX1 U592 ( .IN(Multi_dataout[11]), .OUT(n232) );
  AOI21 U593 ( .IN1(n782), .IN2(n219), .IN3(RSTn_BAR), .OUT(N89) );
  INVX4 U594 ( .IN(n820), .OUT(n482) );
  NANDX2 U595 ( .IN1(n205), .IN2(n482), .OUT(n940) );
  INVX4 U596 ( .IN(n888), .OUT(n746) );
  NANDX2 U597 ( .IN1(n205), .IN2(n746), .OUT(n889) );
  NOR2X1 U598 ( .IN1(n770), .IN2(n769), .OUT(n840) );
  OAI21 U599 ( .IN1(n215), .IN2(n832), .IN3(n839), .OUT(n209) );
  OAI21 U600 ( .IN1(n215), .IN2(N392), .IN3(n218), .OUT(n208) );
  AOI22 U601 ( .IN1(n205), .IN2(n209), .IN3(n745), .IN4(n208), .OUT(n210) );
  OAI21 U602 ( .IN1(n833), .IN2(N392), .IN3(n746), .OUT(n216) );
  INVX4 U603 ( .IN(n219), .OUT(n747) );
  MUX2X1 U604 ( .IN1(n119), .IN2(Final_Exponent_reg[8]), .S(n220), .OUT(n740)
         );
  NOR2X1 U605 ( .IN1(n893), .IN2(Multi_dataout[14]), .OUT(n226) );
  NOR2X1 U606 ( .IN1(Final_Exponent_reg[6]), .IN2(Final_Exponent_reg[7]), 
        .OUT(n228) );
  NOR2X1 U607 ( .IN1(Final_Exponent_reg[4]), .IN2(Final_Exponent_reg[5]), 
        .OUT(n227) );
  NAND3X1 U608 ( .IN1(n119), .IN2(n228), .IN3(n227), .OUT(n229) );
  NOR2X1 U609 ( .IN1(n569), .IN2(n707), .OUT(n647) );
  AOI21 U610 ( .IN1(Final_Exponent_reg[1]), .IN2(n204), .IN3(n413), .OUT(n236)
         );
  NOR2X1 U611 ( .IN1(n486), .IN2(n707), .OUT(n235) );
  NOR2X1 U612 ( .IN1(n236), .IN2(n680), .OUT(n360) );
  OAI21 U613 ( .IN1(Final_Exponent_reg[0]), .IN2(n256), .IN3(n413), .OUT(n401)
         );
  NOR2X1 U614 ( .IN1(Multi_dataout[5]), .IN2(n239), .OUT(n240) );
  AOI21 U615 ( .IN1(n242), .IN2(n103), .IN3(n652), .OUT(n364) );
  NOR2X1 U616 ( .IN1(Multi_dataout[11]), .IN2(n586), .OUT(n243) );
  AOI21 U617 ( .IN1(n416), .IN2(n244), .IN3(n651), .OUT(n385) );
  NOR2X1 U618 ( .IN1(n364), .IN2(n385), .OUT(n253) );
  NOR2X1 U619 ( .IN1(n248), .IN2(n707), .OUT(n654) );
  NOR2X1 U620 ( .IN1(n251), .IN2(n708), .OUT(n658) );
  NAND3X1 U621 ( .IN1(n253), .IN2(n366), .IN3(n387), .OUT(n254) );
  NOR2X1 U622 ( .IN1(Multi_dataout[4]), .IN2(n257), .OUT(n258) );
  NOR2X1 U623 ( .IN1(n435), .IN2(n263), .OUT(n264) );
  NAND3X1 U624 ( .IN1(n268), .IN2(Multi_dataout[0]), .IN3(n447), .OUT(n269) );
  NOR2X1 U625 ( .IN1(n391), .IN2(n57), .OUT(n457) );
  INVX4 U626 ( .IN(n272), .OUT(n379) );
  AOI22 U627 ( .IN1(n598), .IN2(Datain1[10]), .IN3(Datain2[10]), .IN4(n595), 
        .OUT(n286) );
  INVX4 U628 ( .IN(n825), .OUT(n374) );
  NAND3X1 U629 ( .IN1(n277), .IN2(n596), .IN3(n477), .OUT(n620) );
  NOR2X1 U630 ( .IN1(n278), .IN2(n708), .OUT(n279) );
  OAI21 U631 ( .IN1(n281), .IN2(n734), .IN3(n600), .OUT(n282) );
  AOI21 U632 ( .IN1(n622), .IN2(n742), .IN3(n820), .OUT(n283) );
  NOR2X1 U633 ( .IN1(n620), .IN2(n283), .OUT(n294) );
  NAND3X1 U634 ( .IN1(n286), .IN2(n285), .IN3(n284), .OUT(n287) );
  AOI21 U635 ( .IN1(C276_DATA3_3), .IN2(n379), .IN3(n287), .OUT(n288) );
  AOI22 U636 ( .IN1(n351), .IN2(Final_Exponent_reg[3]), .IN3(n205), .IN4(n289), 
        .OUT(n293) );
  INVX4 U637 ( .IN(n380), .OUT(n317) );
  OAI21 U638 ( .IN1(RSTn_BAR), .IN2(n294), .IN3(n895), .OUT(n381) );
  AOI22 U639 ( .IN1(n598), .IN2(DP_OP_357J3_124_4634_n65), .IN3(Datain2[7]), 
        .IN4(n595), .OUT(n297) );
  NAND3X1 U640 ( .IN1(n297), .IN2(n296), .IN3(n295), .OUT(n298) );
  AOI21 U641 ( .IN1(C276_DATA3_0), .IN2(n379), .IN3(n298), .OUT(n299) );
  AOI22 U642 ( .IN1(Final_Exponent_reg[0]), .IN2(n381), .IN3(n205), .IN4(n300), 
        .OUT(n301) );
  AOI22 U643 ( .IN1(n97), .IN2(Final_Exponent_reg[0]), .IN3(
        Final_Exponent_reg[1]), .IN4(n103), .OUT(n303) );
  AOI22 U644 ( .IN1(n598), .IN2(DP_OP_357J3_124_4634_n66), .IN3(
        DP_OP_357J3_124_4634_n58), .IN4(n595), .OUT(n302) );
  OAI21 U645 ( .IN1(n303), .IN2(n332), .IN3(n302), .OUT(n304) );
  AOI21 U646 ( .IN1(N385), .IN2(n374), .IN3(n304), .OUT(n306) );
  AOI22 U647 ( .IN1(Final_Exponent_reg[1]), .IN2(n381), .IN3(n205), .IN4(n307), 
        .OUT(n308) );
  OAI21 U648 ( .IN1(n204), .IN2(n310), .IN3(n309), .OUT(n312) );
  AOI22 U649 ( .IN1(n598), .IN2(Datain1[9]), .IN3(Datain2[9]), .IN4(n595), 
        .OUT(n311) );
  OAI21 U650 ( .IN1(n312), .IN2(n332), .IN3(n311), .OUT(n313) );
  AOI21 U651 ( .IN1(N386), .IN2(n374), .IN3(n313), .OUT(n315) );
  AOI22 U652 ( .IN1(n204), .IN2(n381), .IN3(n205), .IN4(n316), .OUT(n318) );
  AOI22 U653 ( .IN1(n598), .IN2(Datain1[11]), .IN3(Datain2[11]), .IN4(n595), 
        .OUT(n323) );
  OAI21 U654 ( .IN1(n98), .IN2(n319), .IN3(n118), .OUT(n320) );
  NAND3X1 U655 ( .IN1(n321), .IN2(n320), .IN3(n370), .OUT(n322) );
  NAND3X1 U656 ( .IN1(n323), .IN2(n344), .IN3(n322), .OUT(n324) );
  AOI21 U657 ( .IN1(N388), .IN2(n374), .IN3(n324), .OUT(n327) );
  NAND3X1 U658 ( .IN1(n327), .IN2(n326), .IN3(n325), .OUT(n328) );
  AOI22 U659 ( .IN1(n351), .IN2(Final_Exponent_reg[4]), .IN3(n205), .IN4(n328), 
        .OUT(n329) );
  OAI21 U660 ( .IN1(Final_Exponent_reg[5]), .IN2(n330), .IN3(n339), .OUT(n333)
         );
  AOI22 U661 ( .IN1(n598), .IN2(Datain1[12]), .IN3(Datain2[12]), .IN4(n595), 
        .OUT(n331) );
  OAI21 U662 ( .IN1(n333), .IN2(n332), .IN3(n331), .OUT(n334) );
  AOI21 U663 ( .IN1(N389), .IN2(n374), .IN3(n334), .OUT(n335) );
  AOI21 U664 ( .IN1(C276_DATA3_5), .IN2(n379), .IN3(n336), .OUT(n338) );
  AOI21 U665 ( .IN1(Final_Exponent_reg[5]), .IN2(n381), .IN3(n380), .OUT(n337)
         );
  OAI21 U666 ( .IN1(RSTn_BAR), .IN2(n338), .IN3(n337), .OUT(n874) );
  AOI22 U667 ( .IN1(n598), .IN2(Datain1[13]), .IN3(Datain2[13]), .IN4(n595), 
        .OUT(n345) );
  OAI21 U668 ( .IN1(Final_Exponent_reg[6]), .IN2(n342), .IN3(n341), .OUT(n343)
         );
  NAND3X1 U669 ( .IN1(n345), .IN2(n344), .IN3(n343), .OUT(n346) );
  AOI21 U670 ( .IN1(n347), .IN2(Final_Exponent_reg[6]), .IN3(n346), .OUT(n349)
         );
  AOI21 U671 ( .IN1(C276_DATA3_6), .IN2(n379), .IN3(n350), .OUT(n353) );
  OAI21 U672 ( .IN1(RSTn_BAR), .IN2(n353), .IN3(n352), .OUT(n873) );
  NAND3X1 U673 ( .IN1(n361), .IN2(n455), .IN3(n454), .OUT(n354) );
  NAND3X1 U674 ( .IN1(n355), .IN2(n430), .IN3(n357), .OUT(C1_Z_3) );
  NOR2X1 U675 ( .IN1(n450), .IN2(n360), .OUT(n358) );
  NAND3X1 U676 ( .IN1(n358), .IN2(n387), .IN3(n357), .OUT(C1_Z_2) );
  NAND3X1 U677 ( .IN1(n388), .IN2(n384), .IN3(n361), .OUT(n362) );
  NOR2X1 U678 ( .IN1(n368), .IN2(n362), .OUT(n363) );
  NAND3X1 U679 ( .IN1(n366), .IN2(n365), .IN3(n455), .OUT(n367) );
  NOR2X1 U680 ( .IN1(n368), .IN2(n367), .OUT(n369) );
  NAND3X1 U681 ( .IN1(n369), .IN2(n430), .IN3(n429), .OUT(C1_Z_0) );
  AOI22 U682 ( .IN1(n598), .IN2(Datain1[14]), .IN3(Datain2[14]), .IN4(n595), 
        .OUT(n377) );
  MUX2X1 U683 ( .IN1(n373), .IN2(n372), .S(Final_Exponent_reg[7]), .OUT(n376)
         );
  NAND3X1 U684 ( .IN1(n377), .IN2(n376), .IN3(n375), .OUT(n378) );
  AOI21 U685 ( .IN1(C276_DATA3_7), .IN2(n379), .IN3(n378), .OUT(n383) );
  AOI21 U686 ( .IN1(Final_Exponent_reg[7]), .IN2(n381), .IN3(n380), .OUT(n382)
         );
  OAI21 U687 ( .IN1(RSTn_BAR), .IN2(n383), .IN3(n382), .OUT(n872) );
  INVX4 U688 ( .IN(n940), .OUT(n727) );
  NOR2X1 U689 ( .IN1(n386), .IN2(n385), .OUT(n390) );
  NOR2X1 U690 ( .IN1(n392), .IN2(n391), .OUT(n410) );
  NOR2X1 U691 ( .IN1(n393), .IN2(n449), .OUT(n408) );
  AOI21 U692 ( .IN1(n654), .IN2(n395), .IN3(n394), .OUT(n396) );
  AOI21 U693 ( .IN1(n709), .IN2(n401), .IN3(n400), .OUT(n402) );
  NOR2X1 U694 ( .IN1(n403), .IN2(n446), .OUT(n406) );
  OAI21 U695 ( .IN1(n448), .IN2(n692), .IN3(n404), .OUT(n424) );
  NAND3X1 U696 ( .IN1(n406), .IN2(n447), .IN3(n405), .OUT(n407) );
  OAI21 U697 ( .IN1(n408), .IN2(n407), .IN3(Final_Exponent_reg[1]), .OUT(n409)
         );
  OAI21 U698 ( .IN1(n411), .IN2(n648), .IN3(n651), .OUT(n412) );
  NOR2X1 U699 ( .IN1(n412), .IN2(n654), .OUT(n418) );
  NOR2X1 U700 ( .IN1(Final_Exponent_reg[1]), .IN2(n413), .OUT(n415) );
  OAI21 U701 ( .IN1(n416), .IN2(n415), .IN3(n414), .OUT(n417) );
  NOR2X1 U702 ( .IN1(n419), .IN2(n658), .OUT(n423) );
  NAND3X1 U703 ( .IN1(n423), .IN2(n445), .IN3(n422), .OUT(n425) );
  NOR2X1 U704 ( .IN1(n425), .IN2(n424), .OUT(n427) );
  NAND3X1 U705 ( .IN1(n431), .IN2(n430), .IN3(n429), .OUT(n432) );
  AOI21 U706 ( .IN1(Final_Exponent_reg[0]), .IN2(n433), .IN3(n432), .OUT(n441)
         );
  MUX2X1 U707 ( .IN1(n435), .IN2(n434), .S(n439), .OUT(n436) );
  NOR2X1 U708 ( .IN1(n442), .IN2(n436), .OUT(n453) );
  AOI22 U709 ( .IN1(Multi_dataout[2]), .IN2(n605), .IN3(Multi_dataout[5]), 
        .IN4(n521), .OUT(n444) );
  AOI22 U710 ( .IN1(n604), .IN2(Multi_dataout[4]), .IN3(Multi_dataout[3]), 
        .IN4(n603), .OUT(n443) );
  MUX2X1 U711 ( .IN1(n453), .IN2(n518), .S(n488), .OUT(n612) );
  AOI21 U712 ( .IN1(n734), .IN2(Final_Exponent_reg[3]), .IN3(n456), .OUT(n458)
         );
  NOR2X1 U713 ( .IN1(n673), .IN2(n613), .OUT(n463) );
  AOI22 U714 ( .IN1(T_reg), .IN2(n893), .IN3(Multi_dataout[6]), .IN4(n625), 
        .OUT(n460) );
  OAI21 U715 ( .IN1(n461), .IN2(n470), .IN3(n460), .OUT(n462) );
  AOI21 U716 ( .IN1(n612), .IN2(n463), .IN3(n462), .OUT(n696) );
  OAI21 U717 ( .IN1(n712), .IN2(n696), .IN3(n464), .OUT(n124) );
  AOI22 U718 ( .IN1(n604), .IN2(Multi_dataout[1]), .IN3(Multi_dataout[2]), 
        .IN4(n521), .OUT(n465) );
  AOI22 U719 ( .IN1(Multi_dataout[3]), .IN2(n605), .IN3(Multi_dataout[6]), 
        .IN4(n521), .OUT(n468) );
  AOI22 U720 ( .IN1(n604), .IN2(Multi_dataout[5]), .IN3(Multi_dataout[4]), 
        .IN4(n603), .OUT(n467) );
  MUX2X1 U721 ( .IN1(n539), .IN2(n553), .S(n488), .OUT(n473) );
  AOI22 U722 ( .IN1(G_reg), .IN2(n893), .IN3(Multi_dataout[7]), .IN4(n625), 
        .OUT(n469) );
  OAI21 U723 ( .IN1(n471), .IN2(n470), .IN3(n469), .OUT(n472) );
  AOI21 U724 ( .IN1(n473), .IN2(n627), .IN3(n472), .OUT(n697) );
  OAI21 U725 ( .IN1(n712), .IN2(n697), .IN3(n475), .OUT(n125) );
  AOI21 U726 ( .IN1(n476), .IN2(n482), .IN3(n858), .OUT(n478) );
  NAND3X1 U727 ( .IN1(n478), .IN2(n825), .IN3(n477), .OUT(n479) );
  OAI21 U728 ( .IN1(n486), .IN2(n548), .IN3(n485), .OUT(n487) );
  AOI21 U729 ( .IN1(n547), .IN2(Multi_dataout[8]), .IN3(n487), .OUT(n497) );
  AOI22 U730 ( .IN1(Multi_dataout[4]), .IN2(n605), .IN3(Multi_dataout[7]), 
        .IN4(n521), .OUT(n490) );
  AOI22 U731 ( .IN1(n604), .IN2(Multi_dataout[6]), .IN3(Multi_dataout[5]), 
        .IN4(n603), .OUT(n489) );
  INVX4 U732 ( .IN(n492), .OUT(n609) );
  AOI22 U733 ( .IN1(Multi_dataout[0]), .IN2(n605), .IN3(Multi_dataout[3]), 
        .IN4(n521), .OUT(n494) );
  AOI22 U734 ( .IN1(n604), .IN2(Multi_dataout[2]), .IN3(Multi_dataout[1]), 
        .IN4(n603), .OUT(n493) );
  NAND3X1 U735 ( .IN1(n497), .IN2(n496), .IN3(n495), .OUT(n498) );
  AOI22 U736 ( .IN1(Final_Mantissa_reg[0]), .IN2(n618), .IN3(n205), .IN4(n498), 
        .OUT(n499) );
  AOI22 U737 ( .IN1(Multi_dataout[1]), .IN2(n605), .IN3(Multi_dataout[4]), 
        .IN4(n521), .OUT(n501) );
  AOI22 U738 ( .IN1(n604), .IN2(Multi_dataout[3]), .IN3(Multi_dataout[2]), 
        .IN4(n603), .OUT(n500) );
  AOI22 U739 ( .IN1(Multi_dataout[5]), .IN2(n605), .IN3(Multi_dataout[8]), 
        .IN4(n521), .OUT(n503) );
  AOI22 U740 ( .IN1(n604), .IN2(Multi_dataout[7]), .IN3(Multi_dataout[6]), 
        .IN4(n603), .OUT(n502) );
  NAND3X1 U741 ( .IN1(n522), .IN2(n505), .IN3(n744), .OUT(n506) );
  OAI21 U742 ( .IN1(n507), .IN2(n561), .IN3(n506), .OUT(n508) );
  AOI21 U743 ( .IN1(Datain2[1]), .IN2(n595), .IN3(n508), .OUT(n509) );
  OAI21 U744 ( .IN1(n537), .IN2(n548), .IN3(n509), .OUT(n510) );
  AOI21 U745 ( .IN1(n547), .IN2(Multi_dataout[9]), .IN3(n510), .OUT(n511) );
  OAI21 U746 ( .IN1(n512), .IN2(n538), .IN3(n511), .OUT(n513) );
  AOI21 U747 ( .IN1(n611), .IN2(n582), .IN3(n513), .OUT(n514) );
  AOI22 U748 ( .IN1(Final_Mantissa_reg[1]), .IN2(n618), .IN3(n205), .IN4(n516), 
        .OUT(n517) );
  AOI22 U749 ( .IN1(Multi_dataout[6]), .IN2(n605), .IN3(Multi_dataout[9]), 
        .IN4(n521), .OUT(n520) );
  AOI22 U750 ( .IN1(n604), .IN2(Multi_dataout[8]), .IN3(Multi_dataout[7]), 
        .IN4(n603), .OUT(n519) );
  AOI22 U751 ( .IN1(n604), .IN2(Multi_dataout[0]), .IN3(Multi_dataout[1]), 
        .IN4(n521), .OUT(n530) );
  NAND3X1 U752 ( .IN1(n541), .IN2(n523), .IN3(n744), .OUT(n524) );
  OAI21 U753 ( .IN1(n525), .IN2(n561), .IN3(n524), .OUT(n526) );
  AOI21 U754 ( .IN1(Datain2[2]), .IN2(n595), .IN3(n526), .OUT(n527) );
  OAI21 U755 ( .IN1(n569), .IN2(n548), .IN3(n527), .OUT(n528) );
  AOI21 U756 ( .IN1(n547), .IN2(Multi_dataout[10]), .IN3(n528), .OUT(n529) );
  OAI21 U757 ( .IN1(n530), .IN2(n538), .IN3(n529), .OUT(n531) );
  AOI21 U758 ( .IN1(n611), .IN2(n608), .IN3(n531), .OUT(n532) );
  AOI22 U759 ( .IN1(Final_Mantissa_reg[2]), .IN2(n618), .IN3(n205), .IN4(n534), 
        .OUT(n535) );
  AOI22 U760 ( .IN1(n605), .IN2(Multi_dataout[7]), .IN3(Multi_dataout[9]), 
        .IN4(n604), .OUT(n536) );
  OAI21 U761 ( .IN1(n537), .IN2(n585), .IN3(n536), .OUT(n540) );
  AOI22 U762 ( .IN1(n540), .IN2(n611), .IN3(n588), .IN4(n539), .OUT(n555) );
  AOI21 U763 ( .IN1(n541), .IN2(n106), .IN3(n861), .OUT(n543) );
  AOI22 U764 ( .IN1(n543), .IN2(n558), .IN3(Datain1[3]), .IN4(n598), .OUT(n545) );
  AOI21 U765 ( .IN1(n547), .IN2(Multi_dataout[11]), .IN3(n546), .OUT(n551) );
  OAI21 U766 ( .IN1(n581), .IN2(n549), .IN3(n548), .OUT(n602) );
  AOI21 U767 ( .IN1(n609), .IN2(n553), .IN3(n552), .OUT(n554) );
  AOI22 U768 ( .IN1(Final_Mantissa_reg[3]), .IN2(n618), .IN3(n205), .IN4(n556), 
        .OUT(n557) );
  NAND3X1 U769 ( .IN1(n744), .IN2(n577), .IN3(n559), .OUT(n560) );
  OAI21 U770 ( .IN1(n562), .IN2(n561), .IN3(n560), .OUT(n563) );
  AOI21 U771 ( .IN1(Datain2[4]), .IN2(n595), .IN3(n563), .OUT(n564) );
  OAI21 U772 ( .IN1(n58), .IN2(n599), .IN3(n564), .OUT(n566) );
  AOI21 U773 ( .IN1(n602), .IN2(Multi_dataout[11]), .IN3(n566), .OUT(n574) );
  AOI22 U774 ( .IN1(n605), .IN2(Multi_dataout[8]), .IN3(Multi_dataout[10]), 
        .IN4(n604), .OUT(n568) );
  OAI21 U775 ( .IN1(n569), .IN2(n585), .IN3(n568), .OUT(n571) );
  AOI22 U776 ( .IN1(n571), .IN2(n611), .IN3(n588), .IN4(n570), .OUT(n572) );
  NAND3X1 U777 ( .IN1(n574), .IN2(n573), .IN3(n572), .OUT(n575) );
  AOI22 U778 ( .IN1(Final_Mantissa_reg[4]), .IN2(n618), .IN3(n205), .IN4(n575), 
        .OUT(n576) );
  AOI21 U779 ( .IN1(n602), .IN2(n59), .IN3(n579), .OUT(n592) );
  NOR2X1 U780 ( .IN1(n581), .IN2(n580), .OUT(n583) );
  OAI21 U781 ( .IN1(n583), .IN2(n582), .IN3(n609), .OUT(n591) );
  AOI22 U782 ( .IN1(n605), .IN2(Multi_dataout[9]), .IN3(Multi_dataout[11]), 
        .IN4(n604), .OUT(n584) );
  OAI21 U783 ( .IN1(n586), .IN2(n585), .IN3(n584), .OUT(n589) );
  AOI22 U784 ( .IN1(n589), .IN2(n611), .IN3(n588), .IN4(n587), .OUT(n590) );
  NAND3X1 U785 ( .IN1(n592), .IN2(n591), .IN3(n590), .OUT(n593) );
  AOI22 U786 ( .IN1(Final_Mantissa_reg[5]), .IN2(n618), .IN3(n205), .IN4(n593), 
        .OUT(n594) );
  AOI21 U787 ( .IN1(n602), .IN2(Multi_dataout[13]), .IN3(n601), .OUT(n616) );
  AOI22 U788 ( .IN1(n605), .IN2(Multi_dataout[10]), .IN3(Multi_dataout[12]), 
        .IN4(n604), .OUT(n606) );
  AOI22 U789 ( .IN1(n611), .IN2(n610), .IN3(n609), .IN4(n608), .OUT(n615) );
  NAND3X1 U790 ( .IN1(n675), .IN2(n613), .IN3(n612), .OUT(n614) );
  NAND3X1 U791 ( .IN1(n616), .IN2(n615), .IN3(n614), .OUT(n617) );
  AOI22 U792 ( .IN1(Final_Mantissa_reg[6]), .IN2(n618), .IN3(n205), .IN4(n617), 
        .OUT(n619) );
  NAND3X1 U793 ( .IN1(n642), .IN2(n895), .IN3(n621), .OUT(n630) );
  AOI22 U794 ( .IN1(n625), .IN2(n740), .IN3(Final_Exponent_reg[8]), .IN4(n624), 
        .OUT(n629) );
  OAI21 U795 ( .IN1(n825), .IN2(N392), .IN3(n832), .OUT(n635) );
  AOI22 U796 ( .IN1(Exc_value[2]), .IN2(n636), .IN3(n108), .IN4(n635), .OUT(
        n818) );
  OAI21 U797 ( .IN1(n638), .IN2(n835), .IN3(n637), .OUT(n639) );
  AOI21 U798 ( .IN1(n826), .IN2(n120), .IN3(n639), .OUT(n640) );
  OAI21 U799 ( .IN1(n107), .IN2(n810), .IN3(n794), .OUT(ExcCheck_Datain[0]) );
  OAI21 U800 ( .IN1(n111), .IN2(n810), .IN3(n800), .OUT(ExcCheck_Datain[1]) );
  OAI21 U801 ( .IN1(n109), .IN2(n810), .IN3(n801), .OUT(ExcCheck_Datain[2]) );
  OAI21 U802 ( .IN1(n106), .IN2(n810), .IN3(n802), .OUT(ExcCheck_Datain[3]) );
  OAI21 U803 ( .IN1(n112), .IN2(n810), .IN3(n803), .OUT(ExcCheck_Datain[4]) );
  OAI21 U804 ( .IN1(n110), .IN2(n810), .IN3(n804), .OUT(ExcCheck_Datain[5]) );
  OAI21 U805 ( .IN1(n113), .IN2(n810), .IN3(n805), .OUT(ExcCheck_Datain[6]) );
  OAI21 U806 ( .IN1(n103), .IN2(n810), .IN3(n806), .OUT(ExcCheck_Datain[7]) );
  OAI21 U807 ( .IN1(n97), .IN2(n810), .IN3(n807), .OUT(ExcCheck_Datain[8]) );
  OAI21 U808 ( .IN1(n98), .IN2(n810), .IN3(n809), .OUT(ExcCheck_Datain[9]) );
  OAI21 U809 ( .IN1(n102), .IN2(n810), .IN3(n795), .OUT(ExcCheck_Datain[10])
         );
  OAI21 U810 ( .IN1(n118), .IN2(n810), .IN3(n796), .OUT(ExcCheck_Datain[11])
         );
  OAI21 U811 ( .IN1(n116), .IN2(n810), .IN3(n797), .OUT(ExcCheck_Datain[12])
         );
  OAI21 U812 ( .IN1(n100), .IN2(n810), .IN3(n798), .OUT(ExcCheck_Datain[13])
         );
  OAI21 U813 ( .IN1(n117), .IN2(n810), .IN3(n799), .OUT(ExcCheck_Datain[14])
         );
  AOI21 U814 ( .IN1(n745), .IN2(n643), .IN3(n919), .OUT(n641) );
  INVX4 U815 ( .IN(n676), .OUT(n722) );
  AOI21 U816 ( .IN1(n650), .IN2(n719), .IN3(n115), .OUT(n657) );
  AOI21 U817 ( .IN1(n716), .IN2(n657), .IN3(n656), .OUT(n660) );
  AOI22 U818 ( .IN1(n660), .IN2(n720), .IN3(n719), .IN4(n659), .OUT(n661) );
  NOR2X1 U819 ( .IN1(n673), .IN2(n661), .OUT(n662) );
  AOI22 U820 ( .IN1(n115), .IN2(n673), .IN3(n663), .IN4(n662), .OUT(n664) );
  OAI21 U821 ( .IN1(n722), .IN2(n664), .IN3(n695), .OUT(n665) );
  OAI21 U822 ( .IN1(n676), .IN2(n668), .IN3(n666), .OUT(n669) );
  OAI21 U823 ( .IN1(RSOP_428_C1_Z_0), .IN2(n737), .IN3(n669), .OUT(n670) );
  AOI22 U824 ( .IN1(Debug_reg[0]), .IN2(n674), .IN3(n205), .IN4(n670), .OUT(
        n671) );
  AOI22 U825 ( .IN1(Debug_reg[0]), .IN2(n792), .IN3(StateMC[0]), .IN4(n791), 
        .OUT(n672) );
  AOI21 U826 ( .IN1(n678), .IN2(n719), .IN3(n677), .OUT(n701) );
  NAND3X1 U827 ( .IN1(n681), .IN2(n680), .IN3(n679), .OUT(n682) );
  OAI21 U828 ( .IN1(n682), .IN2(n710), .IN3(n719), .OUT(n694) );
  AOI22 U829 ( .IN1(n720), .IN2(n690), .IN3(n719), .IN4(n689), .OUT(n691) );
  OAI21 U830 ( .IN1(n732), .IN2(n692), .IN3(n691), .OUT(n693) );
  AOI22 U831 ( .IN1(Debug_reg[1]), .IN2(n792), .IN3(StateMC[1]), .IN4(n791), 
        .OUT(n704) );
  NOR2X1 U832 ( .IN1(n722), .IN2(Multi_dataout[14]), .OUT(n706) );
  AOI22 U833 ( .IN1(Debug_reg[2]), .IN2(n792), .IN3(StateMC[2]), .IN4(n791), 
        .OUT(n713) );
  NAND3X1 U834 ( .IN1(Debug_reg[3]), .IN2(n715), .IN3(n714), .OUT(n718) );
  NOR2X1 U835 ( .IN1(n718), .IN2(n717), .OUT(n721) );
  AOI22 U836 ( .IN1(n721), .IN2(n720), .IN3(n719), .IN4(n734), .OUT(n724) );
  NAND3X1 U837 ( .IN1(n722), .IN2(Multi_ack), .IN3(Multi_dataout[15]), .OUT(
        n723) );
  OAI21 U838 ( .IN1(n725), .IN2(n724), .IN3(n723), .OUT(n726) );
  AOI22 U839 ( .IN1(Debug_reg[3]), .IN2(n728), .IN3(n727), .IN4(n726), .OUT(
        n729) );
  NOR2X1 U840 ( .IN1(n107), .IN2(n821), .OUT(Dataout[0]) );
  NOR2X1 U841 ( .IN1(n111), .IN2(n821), .OUT(Dataout[1]) );
  NOR2X1 U842 ( .IN1(n109), .IN2(n821), .OUT(Dataout[2]) );
  NOR2X1 U843 ( .IN1(n106), .IN2(n821), .OUT(Dataout[3]) );
  NOR2X1 U844 ( .IN1(n112), .IN2(n821), .OUT(Dataout[4]) );
  NOR2X1 U845 ( .IN1(n110), .IN2(n821), .OUT(Dataout[5]) );
  NOR2X1 U846 ( .IN1(n113), .IN2(n821), .OUT(Dataout[6]) );
  NOR2X1 U847 ( .IN1(n103), .IN2(n821), .OUT(Dataout[7]) );
  NOR2X1 U848 ( .IN1(n97), .IN2(n821), .OUT(Dataout[8]) );
  NOR2X1 U849 ( .IN1(n98), .IN2(n821), .OUT(Dataout[9]) );
  NOR2X1 U850 ( .IN1(n102), .IN2(n821), .OUT(Dataout[10]) );
  NOR2X1 U851 ( .IN1(n118), .IN2(n821), .OUT(Dataout[11]) );
  NOR2X1 U852 ( .IN1(n116), .IN2(n821), .OUT(Dataout[12]) );
  NOR2X1 U853 ( .IN1(n100), .IN2(n821), .OUT(Dataout[13]) );
  NOR2X1 U854 ( .IN1(n117), .IN2(n821), .OUT(Dataout[14]) );
  NOR2X1 U855 ( .IN1(n732), .IN2(n731), .OUT(n733) );
  OAI21 U856 ( .IN1(n171), .IN2(n734), .IN3(n733), .OUT(n735) );
  NAND3X1 U857 ( .IN1(n737), .IN2(n736), .IN3(n735), .OUT(n738) );
  NOR2X1 U858 ( .IN1(n214), .IN2(n215), .OUT(n751) );
  NAND3X1 U859 ( .IN1(Exc_value[0]), .IN2(Exc_value[1]), .IN3(n751), .OUT(n829) );
  INVX1 U860 ( .IN(Exc_value[2]), .OUT(n827) );
  NOR2X1 U861 ( .IN1(n827), .IN2(n213), .OUT(n753) );
  INVX1 U862 ( .IN(Exc_value[0]), .OUT(n836) );
  NAND2X1 U863 ( .IN1(Exc_value[2]), .IN2(n836), .OUT(n752) );
  NOR2X1 U864 ( .IN1(Exc_value[1]), .IN2(n752), .OUT(n854) );
  OAI21 U865 ( .IN1(n829), .IN2(n753), .IN3(n852), .OUT(n856) );
  NAND3X1 U866 ( .IN1(Datain1[10]), .IN2(Datain1[13]), .IN3(Datain1[11]), 
        .OUT(n754) );
  NOR2X1 U867 ( .IN1(n754), .IN2(n765), .OUT(n755) );
  NAND3X1 U868 ( .IN1(DP_OP_357J3_124_4634_n65), .IN2(Datain1[12]), .IN3(n755), 
        .OUT(n763) );
  NOR2X1 U869 ( .IN1(Datain2[9]), .IN2(Datain2[13]), .OUT(n756) );
  NAND3X1 U870 ( .IN1(n758), .IN2(n757), .IN3(n756), .OUT(n762) );
  NOR2X1 U871 ( .IN1(Datain2[14]), .IN2(Datain2[12]), .OUT(n759) );
  NAND3X1 U872 ( .IN1(n759), .IN2(n760), .IN3(n61), .OUT(n761) );
  OAI21 U873 ( .IN1(n60), .IN2(n763), .IN3(n841), .OUT(n777) );
  NOR2X1 U874 ( .IN1(Datain1[13]), .IN2(Datain1[10]), .OUT(n764) );
  NAND3X1 U875 ( .IN1(n60), .IN2(n765), .IN3(n764), .OUT(n770) );
  NOR2X1 U876 ( .IN1(Datain1[14]), .IN2(DP_OP_357J3_124_4634_n65), .OUT(n766)
         );
  NAND3X1 U877 ( .IN1(n767), .IN2(n768), .IN3(n766), .OUT(n769) );
  INVX1 U878 ( .IN(Datain2[14]), .OUT(n775) );
  NAND2X1 U879 ( .IN1(Datain2[10]), .IN2(Datain2[11]), .OUT(n772) );
  NAND3X1 U880 ( .IN1(Datain2[13]), .IN2(DP_OP_357J3_124_4634_n58), .IN3(
        Datain2[9]), .OUT(n771) );
  NOR2X1 U881 ( .IN1(n772), .IN2(n771), .OUT(n773) );
  NAND3X1 U882 ( .IN1(Datain2[12]), .IN2(Datain2[7]), .IN3(n773), .OUT(n774)
         );
  NAND3X1 U883 ( .IN1(n840), .IN2(n775), .IN3(n774), .OUT(n776) );
  OAI21 U884 ( .IN1(Datain1[14]), .IN2(n777), .IN3(n776), .OUT(n833) );
  NAND3X1 U885 ( .IN1(StateMC[1]), .IN2(StateMC[0]), .IN3(n99), .OUT(n891) );
  AOI21 U886 ( .IN1(Multi_dataout[15]), .IN2(n740), .IN3(n893), .OUT(n779) );
  AOI22 U887 ( .IN1(n808), .IN2(n778), .IN3(n890), .IN4(Data_valid), .OUT(n783) );
  OAI21 U888 ( .IN1(n779), .IN2(n894), .IN3(n783), .OUT(n780) );
  NOR2X1 U889 ( .IN1(n781), .IN2(n780), .OUT(n782) );
  AOI21 U890 ( .IN1(n55), .IN2(n784), .IN3(n746), .OUT(n786) );
  AOI22 U891 ( .IN1(n741), .IN2(n740), .IN3(n747), .IN4(n856), .OUT(n785) );
  NAND3X1 U892 ( .IN1(n786), .IN2(n785), .IN3(n820), .OUT(n787) );
  OAI21 U893 ( .IN1(n788), .IN2(n787), .IN3(n205), .OUT(n703) );
  NAND2X1 U894 ( .IN1(Dataout_valid), .IN2(Final_Sign_reg), .OUT(n789) );
  NAND2X1 U895 ( .IN1(Mode[2]), .IN2(n749), .OUT(n790) );
  NOR2X1 U896 ( .IN1(Mode[1]), .IN2(n790), .OUT(n791) );
  AOI21 U897 ( .IN1(Debug_valid_reg), .IN2(n792), .IN3(n791), .OUT(n793) );
  AOI22 U898 ( .IN1(n808), .IN2(Datain1[0]), .IN3(n748), .IN4(Datain2[0]), 
        .OUT(n794) );
  AOI22 U899 ( .IN1(n808), .IN2(Datain1[10]), .IN3(Datain2[10]), .IN4(n748), 
        .OUT(n795) );
  AOI22 U900 ( .IN1(n808), .IN2(Datain1[11]), .IN3(Datain2[11]), .IN4(n748), 
        .OUT(n796) );
  AOI22 U901 ( .IN1(n808), .IN2(Datain1[12]), .IN3(Datain2[12]), .IN4(n748), 
        .OUT(n797) );
  AOI22 U902 ( .IN1(n808), .IN2(Datain1[13]), .IN3(Datain2[13]), .IN4(n748), 
        .OUT(n798) );
  AOI22 U903 ( .IN1(n808), .IN2(Datain1[14]), .IN3(Datain2[14]), .IN4(n748), 
        .OUT(n799) );
  AOI22 U904 ( .IN1(n808), .IN2(Datain1[1]), .IN3(n748), .IN4(Datain2[1]), 
        .OUT(n800) );
  AOI22 U905 ( .IN1(n808), .IN2(Datain1[2]), .IN3(n748), .IN4(Datain2[2]), 
        .OUT(n801) );
  AOI22 U906 ( .IN1(n808), .IN2(Datain1[3]), .IN3(n748), .IN4(Datain2[3]), 
        .OUT(n802) );
  AOI22 U907 ( .IN1(n808), .IN2(Datain1[4]), .IN3(n748), .IN4(Datain2[4]), 
        .OUT(n803) );
  AOI22 U908 ( .IN1(n808), .IN2(Datain1[5]), .IN3(n748), .IN4(Datain2[5]), 
        .OUT(n804) );
  AOI22 U909 ( .IN1(n808), .IN2(Datain1[6]), .IN3(n748), .IN4(Datain2[6]), 
        .OUT(n805) );
  AOI22 U910 ( .IN1(n808), .IN2(DP_OP_357J3_124_4634_n65), .IN3(Datain2[7]), 
        .IN4(n748), .OUT(n806) );
  AOI22 U911 ( .IN1(n808), .IN2(DP_OP_357J3_124_4634_n66), .IN3(
        DP_OP_357J3_124_4634_n58), .IN4(n748), .OUT(n807) );
  AOI22 U912 ( .IN1(n808), .IN2(Datain1[9]), .IN3(Datain2[9]), .IN4(n748), 
        .OUT(n809) );
  NOR2X1 U913 ( .IN1(n215), .IN2(n821), .OUT(Exc[0]) );
  NOR2X1 U914 ( .IN1(n214), .IN2(n821), .OUT(Exc[1]) );
  OAI21 U915 ( .IN1(n850), .IN2(n859), .IN3(n744), .OUT(n811) );
  NOR2X1 U916 ( .IN1(n823), .IN2(n811), .OUT(n838) );
  NOR2X1 U917 ( .IN1(n812), .IN2(n748), .OUT(n813) );
  OAI21 U918 ( .IN1(n55), .IN2(n813), .IN3(n820), .OUT(n822) );
  NOR2X1 U919 ( .IN1(n814), .IN2(n822), .OUT(n832) );
  AOI22 U920 ( .IN1(n213), .IN2(Exc_value[2]), .IN3(n827), .IN4(n108), .OUT(
        n815) );
  NOR2X1 U921 ( .IN1(n829), .IN2(n815), .OUT(n816) );
  NAND3X1 U922 ( .IN1(n818), .IN2(n860), .IN3(n817), .OUT(n819) );
  OAI21 U923 ( .IN1(n838), .IN2(n819), .IN3(n205), .OUT(n667) );
  NAND3X1 U924 ( .IN1(Multi_dataout[15]), .IN2(n742), .IN3(n740), .OUT(n831)
         );
  NOR2X1 U925 ( .IN1(RSTn_BAR), .IN2(n821), .OUT(n830) );
  AOI21 U926 ( .IN1(n823), .IN2(n744), .IN3(n822), .OUT(n824) );
  NAND2X1 U927 ( .IN1(n213), .IN2(n827), .OUT(n828) );
  NOR2X1 U928 ( .IN1(n829), .IN2(n828), .OUT(n853) );
  AOI21 U929 ( .IN1(n747), .IN2(n853), .IN3(Exc[0]), .OUT(n834) );
  OAI21 U930 ( .IN1(n836), .IN2(n835), .IN3(n834), .OUT(n837) );
  NOR2X1 U931 ( .IN1(n838), .IN2(n837), .OUT(n839) );
  NOR2X1 U932 ( .IN1(RSTn_BAR), .IN2(n746), .OUT(n917) );
  AOI21 U933 ( .IN1(n909), .IN2(n841), .IN3(n889), .OUT(n842) );
  AOI21 U934 ( .IN1(Op2_Mantissa_reg[7]), .IN2(n202), .IN3(n842), .OUT(n843)
         );
  OAI21 U935 ( .IN1(Datain2[15]), .IN2(Datain1[15]), .IN3(Data_valid), .OUT(
        n844) );
  AOI21 U936 ( .IN1(Datain2[15]), .IN2(Datain1[15]), .IN3(n844), .OUT(n845) );
  NOR2X1 U937 ( .IN1(RSTn_BAR), .IN2(Data_valid), .OUT(n846) );
  OAI21 U938 ( .IN1(n846), .IN2(n849), .IN3(Final_Sign_reg), .OUT(n847) );
  OAI21 U939 ( .IN1(n849), .IN2(n848), .IN3(n847), .OUT(n880) );
  AOI21 U940 ( .IN1(n854), .IN2(n55), .IN3(n891), .OUT(n858) );
  AOI21 U941 ( .IN1(n55), .IN2(n856), .IN3(n855), .OUT(n857) );
  NOR2X1 U942 ( .IN1(RSTn_BAR), .IN2(n55), .OUT(n887) );
  NAND3X1 U943 ( .IN1(n884), .IN2(n888), .IN3(n861), .OUT(n885) );
  OAI21 U944 ( .IN1(Dataout_valid), .IN2(n885), .IN3(n205), .OUT(n886) );
  MUX2X1 U945 ( .IN1(ExcCheck_valid), .IN2(n887), .S(n886), .OUT(n864) );
  NOR2X1 U946 ( .IN1(StateMC[2]), .IN2(n890), .OUT(n892) );
  AOI21 U947 ( .IN1(n892), .IN2(n891), .IN3(RSTn_BAR), .OUT(n919) );
  OAI21 U948 ( .IN1(n743), .IN2(n939), .IN3(n895), .OUT(n896) );
  NOR2X1 U949 ( .IN1(n920), .IN2(n896), .OUT(n900) );
  AOI21 U950 ( .IN1(n205), .IN2(Multi_ack), .IN3(n896), .OUT(n897) );
  AOI22 U951 ( .IN1(Op1_Mantissa_reg[7]), .IN2(n900), .IN3(Multi_datain1[7]), 
        .IN4(n899), .OUT(n898) );
  AOI22 U952 ( .IN1(n900), .IN2(Op1_Mantissa_reg[6]), .IN3(Multi_datain1[6]), 
        .IN4(n899), .OUT(n901) );
  AOI22 U953 ( .IN1(n745), .IN2(Datain2[6]), .IN3(Op2_Mantissa_reg[6]), .IN4(
        n202), .OUT(n902) );
  AOI22 U954 ( .IN1(n745), .IN2(Datain2[5]), .IN3(Op2_Mantissa_reg[5]), .IN4(
        n202), .OUT(n903) );
  AOI22 U955 ( .IN1(n745), .IN2(Datain2[4]), .IN3(Op2_Mantissa_reg[4]), .IN4(
        n202), .OUT(n904) );
  AOI22 U956 ( .IN1(n745), .IN2(Datain2[3]), .IN3(Op2_Mantissa_reg[3]), .IN4(
        n202), .OUT(n905) );
  AOI22 U957 ( .IN1(n745), .IN2(Datain2[2]), .IN3(Op2_Mantissa_reg[2]), .IN4(
        n202), .OUT(n906) );
  AOI22 U958 ( .IN1(n745), .IN2(Datain2[1]), .IN3(Op2_Mantissa_reg[1]), .IN4(
        n202), .OUT(n907) );
  AOI22 U959 ( .IN1(n745), .IN2(Datain2[0]), .IN3(Op2_Mantissa_reg[0]), .IN4(
        n202), .OUT(n908) );
  AOI22 U960 ( .IN1(n745), .IN2(n909), .IN3(Op1_Mantissa_reg[7]), .IN4(n202), 
        .OUT(n910) );
  AOI22 U961 ( .IN1(n745), .IN2(Datain1[6]), .IN3(Op1_Mantissa_reg[6]), .IN4(
        n202), .OUT(n911) );
  AOI22 U962 ( .IN1(n745), .IN2(Datain1[5]), .IN3(Op1_Mantissa_reg[5]), .IN4(
        n202), .OUT(n912) );
  AOI22 U963 ( .IN1(n745), .IN2(Datain1[4]), .IN3(Op1_Mantissa_reg[4]), .IN4(
        n202), .OUT(n913) );
  AOI22 U964 ( .IN1(n745), .IN2(Datain1[3]), .IN3(Op1_Mantissa_reg[3]), .IN4(
        n202), .OUT(n914) );
  AOI22 U965 ( .IN1(n745), .IN2(Datain1[2]), .IN3(Op1_Mantissa_reg[2]), .IN4(
        n202), .OUT(n915) );
  AOI22 U966 ( .IN1(n745), .IN2(Datain1[1]), .IN3(Op1_Mantissa_reg[1]), .IN4(
        n202), .OUT(n916) );
  AOI22 U967 ( .IN1(n745), .IN2(Datain1[0]), .IN3(Op1_Mantissa_reg[0]), .IN4(
        n202), .OUT(n918) );
  NOR2X1 U968 ( .IN1(n919), .IN2(n745), .OUT(n922) );
  INVX1 U969 ( .IN(n922), .OUT(n921) );
  AOI22 U970 ( .IN1(n922), .IN2(n920), .IN3(Multi_valid_BAR), .IN4(n921), 
        .OUT(n142) );
  NOR2X1 U971 ( .IN1(n921), .IN2(n920), .OUT(n937) );
  OAI21 U972 ( .IN1(RSTn_BAR), .IN2(n750), .IN3(n922), .OUT(n936) );
  AOI22 U973 ( .IN1(Op2_Mantissa_reg[7]), .IN2(n203), .IN3(Multi_datain2[7]), 
        .IN4(n936), .OUT(n923) );
  AOI22 U974 ( .IN1(Op2_Mantissa_reg[6]), .IN2(n203), .IN3(Multi_datain2[6]), 
        .IN4(n936), .OUT(n924) );
  AOI22 U975 ( .IN1(Op2_Mantissa_reg[5]), .IN2(n203), .IN3(Multi_datain2[5]), 
        .IN4(n936), .OUT(n925) );
  AOI22 U976 ( .IN1(Op2_Mantissa_reg[4]), .IN2(n203), .IN3(Multi_datain2[4]), 
        .IN4(n936), .OUT(n926) );
  AOI22 U977 ( .IN1(Op2_Mantissa_reg[3]), .IN2(n203), .IN3(Multi_datain2[3]), 
        .IN4(n936), .OUT(n927) );
  AOI22 U978 ( .IN1(Op2_Mantissa_reg[2]), .IN2(n203), .IN3(Multi_datain2[2]), 
        .IN4(n936), .OUT(n928) );
  AOI22 U979 ( .IN1(Op2_Mantissa_reg[1]), .IN2(n203), .IN3(Multi_datain2[1]), 
        .IN4(n936), .OUT(n929) );
  AOI22 U980 ( .IN1(Op2_Mantissa_reg[0]), .IN2(n203), .IN3(Multi_datain2[0]), 
        .IN4(n936), .OUT(n930) );
  AOI22 U981 ( .IN1(Op1_Mantissa_reg[5]), .IN2(n203), .IN3(Multi_datain1[5]), 
        .IN4(n936), .OUT(n931) );
  AOI22 U982 ( .IN1(Op1_Mantissa_reg[4]), .IN2(n203), .IN3(Multi_datain1[4]), 
        .IN4(n936), .OUT(n932) );
  AOI22 U983 ( .IN1(Op1_Mantissa_reg[3]), .IN2(n203), .IN3(Multi_datain1[3]), 
        .IN4(n936), .OUT(n933) );
  AOI22 U984 ( .IN1(Op1_Mantissa_reg[2]), .IN2(n203), .IN3(Multi_datain1[2]), 
        .IN4(n936), .OUT(n934) );
  AOI22 U985 ( .IN1(Op1_Mantissa_reg[1]), .IN2(n203), .IN3(Multi_datain1[1]), 
        .IN4(n936), .OUT(n935) );
  AOI22 U986 ( .IN1(Op1_Mantissa_reg[0]), .IN2(n203), .IN3(Multi_datain1[0]), 
        .IN4(n936), .OUT(n938) );
endmodule


module FPU_Control ( CLK, RSTn, CS, DIN1, DIN2, DIV, DACK, DR, DOUT, DOV, DOA, 
        ABUSY, MBUSY, EXC, OPT, MODE, DEBUG );
  input [15:0] DIN1;
  input [15:0] DIN2;
  output [15:0] DOUT;
  output [2:0] EXC;
  input [2:0] MODE;
  output [4:0] DEBUG;
  input CLK, RSTn, CS, DIV, DOA, OPT;
  output DACK, DR, DOV, ABUSY, MBUSY;
  wire   Add_carryout, N149, N150, N151, N152, N191, N192, N193,
         MulCntrl_valid, AdderCntrl_valid, AdderCntrl_Dataout_valid,
         MulCntrl_Dataout_valid, Add_valid, Add_ack, AdderCntrl_ExcCheck_valid,
         AdderCntrl_Exc_Ack, Booth_valid, Booth_ack, MulCntrl_ExcCheck_valid,
         MulCntrl_Exc_Ack, ExcSelect, ExcCheck_valid, Booth_Add_valid,
         Booth_Add_ack, AddSelect, u_exc_check_N45, u_exc_check_StateMC_0_,
         u_ExcChecker_interconnect_N53, u_ExcChecker_interconnect_priority_reg,
         u_ExcChecker_interconnect_stateMC_0_,
         u_ExcChecker_interconnect_stateMC_1_, u_booth_N258, u_booth_N55,
         u_booth_N54, u_booth_N53, u_booth_N52, u_booth_N51, u_booth_N50,
         u_booth_N49, u_booth_BStateMC_1_, u_booth_count_reg_2_,
         u_booth_count_reg_3_, u_booth_Q1_reg, u_booth_M_reg_1_,
         u_booth_M_reg_2_, u_booth_M_reg_3_, u_booth_M_reg_4_,
         u_booth_M_reg_5_, u_booth_M_reg_6_, u_booth_M_reg_7_,
         u_booth_A_reg_7_, u_booth_A_reg_8_, u_adder_24b_N131,
         u_adder_24b_N130, u_adder_24b_N129, u_adder_24b_N128,
         u_adder_24b_N127, u_adder_24b_N126, u_adder_24b_N125,
         u_adder_24b_N124, u_adder_24b_N123, u_adder_24b_N122, u_adder_24b_N52,
         u_adder_24b_StateMC_1_, u_Adder_interconnect_N53,
         u_Adder_interconnect_priority_reg, u_Adder_interconnect_stateMC_1_,
         n408, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n462, n463,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n587, n588, n592, n594,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n610,
         n611, n612, n613, n614, n615, n616, n617, n622, n654, n694, n695,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n732, n768, n802, n806, n992, n1022,
         n1028, n1031, n1034, n1037, n1040, n1043, n1077, n1079, n1088, n1092,
         n1135, n1302, n1513, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1587, n1588, n1589, n1620,
         n1621, n1622, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1692, n1723, add_x_176_n13, add_x_176_n12, add_x_176_n11,
         add_x_176_n10, add_x_176_n9, add_x_176_n8, add_x_176_n7, add_x_176_n6,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2;
  wire   [8:0] Add_dataout;
  wire   [4:0] AdderCntrl_Debug;
  wire   [1:0] multStateMC;
  wire   [4:0] MulCntrl_Debug;
  wire   [15:0] AdderCntrl_Op1;
  wire   [15:0] AdderCntrl_Op2;
  wire   [15:0] MulCntrl_Op1;
  wire   [15:0] MulCntrl_Op2;
  wire   [1:0] getdataStat_reg;
  wire   [15:0] AdderResult_reg;
  wire   [15:0] MultResult_reg;
  wire   [2:0] AddExc_reg;
  wire   [2:0] MultExc_reg;
  wire   [15:0] AdderCntrl_Dataout;
  wire   [2:0] AdderCntrl_Exc;
  wire   [15:0] MulCntrl_Dataout;
  wire   [2:0] MulCntrl_Exc;
  wire   [7:0] Add_Op1;
  wire   [8:0] Add_Op2;
  wire   [14:0] AdderCntrl_ExcCheck_Datain;
  wire   [2:0] ExcCheck_value;
  wire   [7:0] Booth_datain1;
  wire   [7:0] Booth_datain2;
  wire   [15:0] Booth_dataout;
  wire   [14:0] MulCntrl_ExcCheck_Datain;
  wire   [8:1] Booth_Add_datain1;
  wire   [8:1] Booth_Add_datain2;
  wire   [8:0] Add_Op1_wire;
  wire   [8:0] Add_Op2_wire;

  Adder_cntrl u_adder_cntrl ( .CLK(CLK), .Datain1({AdderCntrl_Op1[15:13], 
        n1742, AdderCntrl_Op1[11], n1744, n1746, n1810, n1808, 
        AdderCntrl_Op1[6:0]}), .Datain2({AdderCntrl_Op2[15:12], n1739, n1740, 
        AdderCntrl_Op2[9], n1809, n1815, AdderCntrl_Op2[6:0]}), .Data_valid(
        AdderCntrl_valid), .Dataout(AdderCntrl_Dataout), .Dataout_valid(
        AdderCntrl_Dataout_valid), .Exc(AdderCntrl_Exc), .Mode(MODE), .Debug(
        AdderCntrl_Debug), .Adder_datain1({SYNOPSYS_UNCONNECTED_1, Add_Op1}), 
        .Adder_datain2(Add_Op2), .Adder_valid(Add_valid), .Adder_dataout(
        Add_dataout), .Adder_carryout(Add_carryout), .Adder_ack(Add_ack), 
        .ExcCheck_valid(AdderCntrl_ExcCheck_valid), .Exc_value(ExcCheck_value), 
        .Exc_Ack(AdderCntrl_Exc_Ack), .RSTn_BAR(n1833), .ExcCheck_Datain_14_(
        AdderCntrl_ExcCheck_Datain[14]), .ExcCheck_Datain_13__BAR(
        AdderCntrl_ExcCheck_Datain[13]), .ExcCheck_Datain_12_(
        AdderCntrl_ExcCheck_Datain[12]), .ExcCheck_Datain_11_(
        AdderCntrl_ExcCheck_Datain[11]), .ExcCheck_Datain_9_(
        AdderCntrl_ExcCheck_Datain[9]), .ExcCheck_Datain_8_(
        AdderCntrl_ExcCheck_Datain[8]), .ExcCheck_Datain_6_(
        AdderCntrl_ExcCheck_Datain[6]), .ExcCheck_Datain_5_(
        AdderCntrl_ExcCheck_Datain[5]), .ExcCheck_Datain_4_(
        AdderCntrl_ExcCheck_Datain[4]), .ExcCheck_Datain_3_(
        AdderCntrl_ExcCheck_Datain[3]), .ExcCheck_Datain_2_(
        AdderCntrl_ExcCheck_Datain[2]), .ExcCheck_Datain_1_(
        AdderCntrl_ExcCheck_Datain[1]), .ExcCheck_Datain_0_(
        AdderCntrl_ExcCheck_Datain[0]), .ExcCheck_Datain_10__BAR(
        AdderCntrl_ExcCheck_Datain[10]), .ExcCheck_Datain_7__BAR(
        AdderCntrl_ExcCheck_Datain[7]) );
  Mul_cntrl u_mul_cntrl ( .CLK(CLK), .Datain1({MulCntrl_Op1[15:14], n1814, 
        n1817, n1812, MulCntrl_Op1[10:0]}), .Datain2({MulCntrl_Op2[15:13], 
        n1738, n1737, n1734, n1735, MulCntrl_Op2[8], n1818, MulCntrl_Op2[6:0]}), .Data_valid(MulCntrl_valid), .Dataout(MulCntrl_Dataout), .Dataout_valid(
        MulCntrl_Dataout_valid), .Exc(MulCntrl_Exc), .Mode(MODE), .Debug(
        MulCntrl_Debug), .Multi_datain1(Booth_datain1), .Multi_datain2(
        Booth_datain2), .Multi_dataout(Booth_dataout), .Multi_ack(Booth_ack), 
        .ExcCheck_valid(MulCntrl_ExcCheck_valid), .ExcCheck_Datain({
        SYNOPSYS_UNCONNECTED_2, MulCntrl_ExcCheck_Datain}), .Exc_value(
        ExcCheck_value), .RSTn_BAR(n1833), .Multi_valid_BAR(Booth_valid), 
        .Exc_Ack_BAR(n1730) );
  DFFRX1 u_Adder_interconnect_M2_ack_reg ( .D(n1587), .CLK(CLK), .CLRB(n408), 
        .Q(Booth_Add_ack), .QB(n1766) );
  DFFRX1 u_booth_count_reg_reg_0_ ( .D(n1554), .CLK(CLK), .CLRB(n408), .QB(
        n694) );
  DFFRX1 u_booth_count_reg_reg_1_ ( .D(n1079), .CLK(CLK), .CLRB(n408), .Q(n695) );
  DFFRX1 u_booth_count_reg_reg_2_ ( .D(n1555), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_count_reg_2_) );
  DFFRX1 u_booth_count_reg_reg_3_ ( .D(n1092), .CLK(CLK), .CLRB(n408), .Q(
        n1789), .QB(u_booth_count_reg_3_) );
  DFFRX1 u_booth_BStateMC_reg_0_ ( .D(n1556), .CLK(CLK), .CLRB(n408), .Q(n1765), .QB(n732) );
  DFFRX1 u_booth_BStateMC_reg_1_ ( .D(n1088), .CLK(CLK), .CLRB(n408), .Q(n1779), .QB(u_booth_BStateMC_1_) );
  DFFRX1 u_booth_Q_reg_reg_7_ ( .D(n1022), .CLK(CLK), .CLRB(n408), .Q(n720), 
        .QB(n1781) );
  DFFRX1 u_booth_Q_reg_reg_6_ ( .D(n1028), .CLK(CLK), .CLRB(n408), .Q(n719), 
        .QB(n1782) );
  DFFRX1 u_booth_Q_reg_reg_5_ ( .D(n1031), .CLK(CLK), .CLRB(n408), .Q(n718), 
        .QB(n1783) );
  DFFRX1 u_booth_Q_reg_reg_4_ ( .D(n1034), .CLK(CLK), .CLRB(n408), .Q(n717), 
        .QB(n1784) );
  DFFRX1 u_booth_Q_reg_reg_3_ ( .D(n1037), .CLK(CLK), .CLRB(n408), .Q(n716), 
        .QB(n1785) );
  DFFRX1 u_booth_Q_reg_reg_2_ ( .D(n1040), .CLK(CLK), .CLRB(n408), .Q(n715), 
        .QB(n1786) );
  DFFRX1 u_booth_Q_reg_reg_1_ ( .D(n1043), .CLK(CLK), .CLRB(n408), .Q(n714), 
        .QB(n1787) );
  DFFRX1 u_booth_Q_reg_reg_0_ ( .D(n1135), .CLK(CLK), .CLRB(n408), .Q(n713), 
        .QB(n1753) );
  DFFRX1 u_booth_Adder_valid_reg ( .D(n1653), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_valid), .QB(n1780) );
  DFFRX1 u_Adder_interconnect_priority_reg_reg ( .D(n1620), .CLK(CLK), .CLRB(
        n408), .Q(u_Adder_interconnect_priority_reg), .QB(n1757) );
  DFFRX1 u_Adder_interconnect_stateMC_reg_0_ ( .D(n1621), .CLK(CLK), .CLRB(
        n408), .Q(n1756), .QB(n806) );
  DFFRX1 u_Adder_interconnect_M1_ack_reg ( .D(n594), .CLK(CLK), .CLRB(n408), 
        .Q(Add_ack) );
  DFFRX1 u_ExcChecker_interconnect_stateMC_reg_1_ ( .D(n1661), .CLK(CLK), 
        .CLRB(n408), .Q(u_ExcChecker_interconnect_stateMC_1_), .QB(n1775) );
  DFFRX1 u_ExcChecker_interconnect_priority_reg_reg ( .D(n1659), .CLK(CLK), 
        .CLRB(n408), .Q(u_ExcChecker_interconnect_priority_reg), .QB(n1772) );
  DFFRX1 u_ExcChecker_interconnect_stateMC_reg_0_ ( .D(n1660), .CLK(CLK), 
        .CLRB(n408), .Q(u_ExcChecker_interconnect_stateMC_0_), .QB(n1773) );
  DFFRX1 u_ExcChecker_interconnect_S_req_reg ( .D(
        u_ExcChecker_interconnect_N53), .CLK(CLK), .CLRB(n408), .Q(
        ExcCheck_valid) );
  DFFRX1 u_exc_check_ACK_reg ( .D(u_exc_check_N45), .CLK(CLK), .CLRB(n408), 
        .QB(n1769) );
  DFFRX1 u_ExcChecker_interconnect_M2_ack_reg ( .D(n1656), .CLK(CLK), .CLRB(
        n408), .Q(MulCntrl_Exc_Ack), .QB(n1730) );
  DFFRX1 u_exc_check_StateMC_reg_0_ ( .D(n622), .CLK(CLK), .CLRB(n408), .Q(
        u_exc_check_StateMC_0_), .QB(n1788) );
  DFFRX1 u_exc_check_StateMC_reg_1_ ( .D(n1657), .CLK(CLK), .CLRB(n408), .Q(
        n1794), .QB(n654) );
  DFFRX1 u_ExcChecker_interconnect_Select_reg ( .D(n1658), .CLK(CLK), .CLRB(
        n408), .Q(ExcSelect), .QB(n1768) );
  DFFRX1 u_exc_check_AEXC_reg_2_ ( .D(n588), .CLK(CLK), .CLRB(n408), .Q(
        ExcCheck_value[2]) );
  DFFRX1 u_exc_check_AEXC_reg_1_ ( .D(n1654), .CLK(CLK), .CLRB(n408), .Q(
        ExcCheck_value[1]), .QB(n1778) );
  DFFRX1 u_exc_check_AEXC_reg_0_ ( .D(n1655), .CLK(CLK), .CLRB(n408), .Q(
        ExcCheck_value[0]), .QB(n1791) );
  DFFRX1 u_ExcChecker_interconnect_M1_ack_reg ( .D(n592), .CLK(CLK), .CLRB(
        n408), .Q(AdderCntrl_Exc_Ack) );
  DFFRX1 u_Adder_interconnect_stateMC_reg_1_ ( .D(n1622), .CLK(CLK), .CLRB(
        n408), .Q(u_Adder_interconnect_stateMC_1_), .QB(n1774) );
  DFFRX1 u_Adder_interconnect_S_req_reg ( .D(u_Adder_interconnect_N53), .CLK(
        CLK), .CLRB(n408), .Q(n1759), .QB(n802) );
  DFFRX1 u_adder_24b_StateMC_reg_1_ ( .D(n1589), .CLK(CLK), .CLRB(n408), .Q(
        u_adder_24b_StateMC_1_), .QB(n1777) );
  DFFRX1 u_adder_24b_StateMC_reg_0_ ( .D(n1588), .CLK(CLK), .CLRB(n408), .Q(
        n1792), .QB(n768) );
  DFFRX1 u_adder_24b_ACK_reg ( .D(u_adder_24b_N52), .CLK(CLK), .CLRB(n408), 
        .QB(n1770) );
  DFFRX1 u_adder_24b_Z_reg_8_ ( .D(n598), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[8]) );
  DFFRX1 u_adder_24b_Z_reg_7_ ( .D(n599), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[7]) );
  DFFRX1 u_adder_24b_Z_reg_6_ ( .D(n600), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[6]) );
  DFFRX1 u_adder_24b_Z_reg_5_ ( .D(n601), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[5]) );
  DFFRX1 u_adder_24b_Z_reg_4_ ( .D(n602), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[4]) );
  DFFRX1 u_adder_24b_Z_reg_3_ ( .D(n603), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[3]) );
  DFFRX1 u_adder_24b_Z_reg_2_ ( .D(n604), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[2]) );
  DFFRX1 u_adder_24b_Z_reg_1_ ( .D(n605), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[1]) );
  DFFRX1 u_adder_24b_Z_reg_0_ ( .D(n596), .CLK(CLK), .CLRB(n408), .Q(
        Add_dataout[0]) );
  DFFRX1 u_adder_24b_COUT_reg ( .D(n597), .CLK(CLK), .CLRB(n408), .Q(
        Add_carryout) );
  DFFRX1 adderStateMC_reg_0_ ( .D(n1302), .CLK(CLK), .CLRB(n408), .Q(n463), 
        .QB(n1764) );
  DFFRX1 outputRdy_reg_reg_0_ ( .D(N191), .CLK(CLK), .CLRB(n408), .QB(n587) );
  DFFRX1 adderStateMC_reg_1_ ( .D(n1692), .CLK(CLK), .CLRB(n408), .Q(n1761), 
        .QB(n462) );
  DFFRX1 getdataStat_reg_reg_0_ ( .D(N149), .CLK(CLK), .CLRB(n408), .Q(
        getdataStat_reg[0]) );
  DFFRX1 AdderCntrl_Op2_reg_0_ ( .D(n551), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[0]) );
  DFFRX1 AdderCntrl_Op2_reg_1_ ( .D(n550), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[1]) );
  DFFRX1 AdderCntrl_Op2_reg_2_ ( .D(n549), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[2]) );
  DFFRX1 AdderCntrl_Op2_reg_3_ ( .D(n548), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[3]) );
  DFFRX1 AdderCntrl_Op2_reg_4_ ( .D(n547), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[4]) );
  DFFRX1 AdderCntrl_Op2_reg_5_ ( .D(n546), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[5]) );
  DFFRX1 AdderCntrl_Op2_reg_6_ ( .D(n545), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[6]) );
  DFFRX1 AdderCntrl_Op2_reg_7_ ( .D(n544), .CLK(CLK), .CLRB(n408), .QB(n1752)
         );
  DFFRX1 AdderCntrl_Op2_reg_8_ ( .D(n543), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[8]) );
  DFFRX1 AdderCntrl_Op2_reg_9_ ( .D(n542), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[9]) );
  DFFRX1 AdderCntrl_Op2_reg_10_ ( .D(n541), .CLK(CLK), .CLRB(n408), .QB(n1733)
         );
  DFFRX1 AdderCntrl_Op2_reg_11_ ( .D(n540), .CLK(CLK), .CLRB(n408), .QB(n1736)
         );
  DFFRX1 AdderCntrl_Op2_reg_12_ ( .D(n539), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[12]) );
  DFFRX1 AdderCntrl_Op2_reg_13_ ( .D(n538), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[13]) );
  DFFRX1 AdderCntrl_Op2_reg_14_ ( .D(n537), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[14]) );
  DFFRX1 AdderCntrl_Op2_reg_15_ ( .D(n536), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op2[15]) );
  DFFRX1 AdderCntrl_Op1_reg_0_ ( .D(n535), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[0]) );
  DFFRX1 AdderCntrl_Op1_reg_1_ ( .D(n534), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[1]) );
  DFFRX1 AdderCntrl_Op1_reg_2_ ( .D(n533), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[2]) );
  DFFRX1 AdderCntrl_Op1_reg_3_ ( .D(n532), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[3]) );
  DFFRX1 AdderCntrl_Op1_reg_4_ ( .D(n531), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[4]) );
  DFFRX1 AdderCntrl_Op1_reg_5_ ( .D(n530), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[5]) );
  DFFRX1 AdderCntrl_Op1_reg_6_ ( .D(n529), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[6]) );
  DFFRX1 AdderCntrl_Op1_reg_7_ ( .D(n528), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[7]) );
  DFFRX1 AdderCntrl_Op1_reg_8_ ( .D(n527), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[8]) );
  DFFRX1 AdderCntrl_Op1_reg_9_ ( .D(n526), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[9]), .QB(n1745) );
  DFFRX1 AdderCntrl_Op1_reg_10_ ( .D(n525), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[10]), .QB(n1743) );
  DFFRX1 AdderCntrl_Op1_reg_11_ ( .D(n524), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[11]) );
  DFFRX1 AdderCntrl_Op1_reg_12_ ( .D(n523), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[12]), .QB(n1741) );
  DFFRX1 AdderCntrl_Op1_reg_13_ ( .D(n522), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[13]) );
  DFFRX1 AdderCntrl_Op1_reg_14_ ( .D(n521), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[14]) );
  DFFRX1 AdderCntrl_Op1_reg_15_ ( .D(n520), .CLK(CLK), .CLRB(n408), .Q(
        AdderCntrl_Op1[15]) );
  DFFRX1 ABUSY_reg ( .D(N151), .CLK(CLK), .CLRB(n408), .Q(ABUSY) );
  DFFRX1 AddExc_reg_reg_2_ ( .D(n414), .CLK(CLK), .CLRB(n408), .Q(
        AddExc_reg[2]) );
  DFFRX1 AddExc_reg_reg_1_ ( .D(n413), .CLK(CLK), .CLRB(n408), .Q(
        AddExc_reg[1]) );
  DFFRX1 AddExc_reg_reg_0_ ( .D(n412), .CLK(CLK), .CLRB(n408), .Q(
        AddExc_reg[0]) );
  DFFRX1 AdderResult_reg_reg_0_ ( .D(n415), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[0]) );
  DFFRX1 AdderResult_reg_reg_1_ ( .D(n416), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[1]) );
  DFFRX1 AdderResult_reg_reg_2_ ( .D(n417), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[2]) );
  DFFRX1 AdderResult_reg_reg_3_ ( .D(n418), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[3]) );
  DFFRX1 AdderResult_reg_reg_4_ ( .D(n419), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[4]) );
  DFFRX1 AdderResult_reg_reg_5_ ( .D(n420), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[5]) );
  DFFRX1 AdderResult_reg_reg_6_ ( .D(n421), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[6]) );
  DFFRX1 AdderResult_reg_reg_7_ ( .D(n422), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[7]) );
  DFFRX1 AdderResult_reg_reg_8_ ( .D(n423), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[8]) );
  DFFRX1 AdderResult_reg_reg_9_ ( .D(n424), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[9]) );
  DFFRX1 AdderResult_reg_reg_10_ ( .D(n425), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[10]) );
  DFFRX1 AdderResult_reg_reg_11_ ( .D(n426), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[11]) );
  DFFRX1 AdderResult_reg_reg_12_ ( .D(n427), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[12]) );
  DFFRX1 AdderResult_reg_reg_13_ ( .D(n428), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[13]) );
  DFFRX1 AdderResult_reg_reg_14_ ( .D(n429), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[14]) );
  DFFRX1 AdderResult_reg_reg_15_ ( .D(n430), .CLK(CLK), .CLRB(n408), .Q(
        AdderResult_reg[15]) );
  DFFRX1 u_booth_Q1_reg_reg ( .D(n1077), .CLK(CLK), .CLRB(n408), .Q(n1763), 
        .QB(u_booth_Q1_reg) );
  DFFRX1 u_booth_A_reg_reg_8_ ( .D(n1545), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_A_reg_8_), .QB(n1793) );
  DFFRX1 u_booth_A_reg_reg_7_ ( .D(n1546), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_A_reg_7_), .QB(n1776) );
  DFFRX1 u_booth_A_reg_reg_6_ ( .D(n1547), .CLK(CLK), .CLRB(n408), .Q(n1796), 
        .QB(n728) );
  DFFRX1 u_booth_A_reg_reg_5_ ( .D(n1548), .CLK(CLK), .CLRB(n408), .Q(n1795), 
        .QB(n727) );
  DFFRX1 u_booth_A_reg_reg_4_ ( .D(n1549), .CLK(CLK), .CLRB(n408), .Q(n1800), 
        .QB(n726) );
  DFFRX1 u_booth_A_reg_reg_3_ ( .D(n1550), .CLK(CLK), .CLRB(n408), .Q(n1797), 
        .QB(n725) );
  DFFRX1 u_booth_A_reg_reg_2_ ( .D(n1551), .CLK(CLK), .CLRB(n408), .Q(n1798), 
        .QB(n724) );
  DFFRX1 u_booth_A_reg_reg_1_ ( .D(n1552), .CLK(CLK), .CLRB(n408), .Q(n1799), 
        .QB(n723) );
  DFFRX1 u_booth_A_reg_reg_0_ ( .D(n1553), .CLK(CLK), .CLRB(n408), .Q(n1801), 
        .QB(n722) );
  DFFRX1 u_booth_Adder_datain1_reg_0_ ( .D(u_booth_N49), .CLK(CLK), .CLRB(n408), .QB(n1758) );
  DFFRX1 u_booth_Q_reg_reg_8_ ( .D(n1544), .CLK(CLK), .CLRB(n408), .Q(n1790), 
        .QB(n721) );
  DFFRX1 u_booth_Adder_datain1_reg_1_ ( .D(u_booth_N50), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[1]) );
  DFFRX1 u_booth_Adder_datain1_reg_2_ ( .D(u_booth_N51), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[2]) );
  DFFRX1 u_booth_Adder_datain1_reg_3_ ( .D(u_booth_N52), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[3]) );
  DFFRX1 u_booth_Adder_datain1_reg_4_ ( .D(u_booth_N53), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[4]) );
  DFFRX1 u_booth_Adder_datain1_reg_5_ ( .D(u_booth_N54), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[5]) );
  DFFRX1 u_booth_Adder_datain1_reg_6_ ( .D(u_booth_N55), .CLK(CLK), .CLRB(n408), .Q(Booth_Add_datain1[6]) );
  DFFRX1 u_booth_Adder_datain1_reg_7_ ( .D(n706), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain1[7]) );
  DFFRX1 u_booth_Adder_datain1_reg_8_ ( .D(n707), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain1[8]) );
  DFFRX1 u_booth_Adder_datain2_reg_8_ ( .D(n705), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[8]) );
  DFFRX1 u_booth_M_reg_reg_0_ ( .D(n610), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_N258), .QB(n1754) );
  DFFRX1 u_booth_Adder_datain2_reg_0_ ( .D(n697), .CLK(CLK), .CLRB(n408), .QB(
        n1760) );
  DFFRX1 u_booth_M_reg_reg_1_ ( .D(n611), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_1_), .QB(n1762) );
  DFFRX1 u_booth_Adder_datain2_reg_1_ ( .D(n698), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[1]) );
  DFFRX1 u_booth_M_reg_reg_2_ ( .D(n612), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_2_) );
  DFFRX1 u_booth_Adder_datain2_reg_2_ ( .D(n699), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[2]) );
  DFFRX1 u_booth_M_reg_reg_3_ ( .D(n613), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_3_) );
  DFFRX1 u_booth_Adder_datain2_reg_3_ ( .D(n700), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[3]) );
  DFFRX1 u_booth_M_reg_reg_4_ ( .D(n614), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_4_) );
  DFFRX1 u_booth_Adder_datain2_reg_4_ ( .D(n701), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[4]) );
  DFFRX1 u_booth_M_reg_reg_5_ ( .D(n615), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_5_) );
  DFFRX1 u_booth_Adder_datain2_reg_5_ ( .D(n702), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[5]) );
  DFFRX1 u_booth_M_reg_reg_6_ ( .D(n616), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_6_) );
  DFFRX1 u_booth_Adder_datain2_reg_6_ ( .D(n703), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[6]) );
  DFFRX1 u_booth_M_reg_reg_7_ ( .D(n617), .CLK(CLK), .CLRB(n408), .Q(
        u_booth_M_reg_7_), .QB(n1771) );
  DFFRX1 u_booth_Adder_datain2_reg_7_ ( .D(n704), .CLK(CLK), .CLRB(n408), .Q(
        Booth_Add_datain2[7]) );
  DFFRX1 multStateMC_reg_0_ ( .D(n992), .CLK(CLK), .CLRB(n408), .Q(n1767), 
        .QB(multStateMC[0]) );
  DFFRX1 outputRdy_reg_reg_1_ ( .D(N192), .CLK(CLK), .CLRB(n408), .QB(n584) );
  DFFRX1 multStateMC_reg_1_ ( .D(n1513), .CLK(CLK), .CLRB(n408), .Q(
        multStateMC[1]), .QB(n1755) );
  DFFRX1 getdataStat_reg_reg_1_ ( .D(N150), .CLK(CLK), .CLRB(n408), .Q(
        getdataStat_reg[1]) );
  DFFRX1 MulCntrl_Op2_reg_0_ ( .D(n583), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[0]) );
  DFFRX1 MulCntrl_Op2_reg_1_ ( .D(n582), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[1]) );
  DFFRX1 MulCntrl_Op2_reg_2_ ( .D(n581), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[2]) );
  DFFRX1 MulCntrl_Op2_reg_3_ ( .D(n580), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[3]) );
  DFFRX1 MulCntrl_Op2_reg_4_ ( .D(n579), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[4]) );
  DFFRX1 MulCntrl_Op2_reg_5_ ( .D(n578), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[5]) );
  DFFRX1 MulCntrl_Op2_reg_6_ ( .D(n577), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[6]) );
  DFFRX1 MulCntrl_Op2_reg_7_ ( .D(n576), .CLK(CLK), .CLRB(n408), .QB(n1751) );
  DFFRX1 MulCntrl_Op2_reg_8_ ( .D(n575), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[8]) );
  DFFRX1 MulCntrl_Op2_reg_9_ ( .D(n574), .CLK(CLK), .CLRB(n408), .Q(n1735) );
  DFFRX1 MulCntrl_Op2_reg_10_ ( .D(n573), .CLK(CLK), .CLRB(n408), .Q(n1734) );
  DFFRX1 MulCntrl_Op2_reg_11_ ( .D(n572), .CLK(CLK), .CLRB(n408), .Q(n1737) );
  DFFRX1 MulCntrl_Op2_reg_12_ ( .D(n571), .CLK(CLK), .CLRB(n408), .Q(n1738) );
  DFFRX1 MulCntrl_Op2_reg_13_ ( .D(n570), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[13]) );
  DFFRX1 MulCntrl_Op2_reg_14_ ( .D(n569), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[14]) );
  DFFRX1 MulCntrl_Op2_reg_15_ ( .D(n568), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op2[15]) );
  DFFRX1 MulCntrl_Op1_reg_0_ ( .D(n567), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[0]) );
  DFFRX1 MulCntrl_Op1_reg_1_ ( .D(n566), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[1]) );
  DFFRX1 MulCntrl_Op1_reg_2_ ( .D(n565), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[2]) );
  DFFRX1 MulCntrl_Op1_reg_3_ ( .D(n564), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[3]) );
  DFFRX1 MulCntrl_Op1_reg_4_ ( .D(n563), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[4]) );
  DFFRX1 MulCntrl_Op1_reg_5_ ( .D(n562), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[5]) );
  DFFRX1 MulCntrl_Op1_reg_6_ ( .D(n561), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[6]) );
  DFFRX1 MulCntrl_Op1_reg_7_ ( .D(n560), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[7]) );
  DFFRX1 MulCntrl_Op1_reg_8_ ( .D(n559), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[8]) );
  DFFRX1 MulCntrl_Op1_reg_9_ ( .D(n558), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[9]) );
  DFFRX1 MulCntrl_Op1_reg_10_ ( .D(n557), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[10]) );
  DFFRX1 MulCntrl_Op1_reg_11_ ( .D(n556), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[11]), .QB(n1811) );
  DFFRX1 MulCntrl_Op1_reg_12_ ( .D(n555), .CLK(CLK), .CLRB(n408), .QB(n1813)
         );
  DFFRX1 MulCntrl_Op1_reg_13_ ( .D(n554), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[13]) );
  DFFRX1 MulCntrl_Op1_reg_14_ ( .D(n553), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[14]) );
  DFFRX1 MulCntrl_Op1_reg_15_ ( .D(n552), .CLK(CLK), .CLRB(n408), .Q(
        MulCntrl_Op1[15]) );
  DFFRX1 MBUSY_reg ( .D(N152), .CLK(CLK), .CLRB(n408), .Q(MBUSY) );
  DFFRX1 DR_reg ( .D(N193), .CLK(CLK), .CLRB(n408), .Q(DR) );
  DFFRX1 MultExc_reg_reg_2_ ( .D(n469), .CLK(CLK), .CLRB(n408), .Q(
        MultExc_reg[2]) );
  DFFRX1 MultExc_reg_reg_1_ ( .D(n468), .CLK(CLK), .CLRB(n408), .Q(
        MultExc_reg[1]) );
  DFFRX1 MultExc_reg_reg_0_ ( .D(n467), .CLK(CLK), .CLRB(n408), .Q(
        MultExc_reg[0]) );
  DFFRX1 MultResult_reg_reg_0_ ( .D(n470), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[0]) );
  DFFRX1 MultResult_reg_reg_1_ ( .D(n471), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[1]) );
  DFFRX1 MultResult_reg_reg_2_ ( .D(n472), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[2]) );
  DFFRX1 MultResult_reg_reg_3_ ( .D(n473), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[3]) );
  DFFRX1 MultResult_reg_reg_4_ ( .D(n474), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[4]) );
  DFFRX1 MultResult_reg_reg_5_ ( .D(n475), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[5]) );
  DFFRX1 MultResult_reg_reg_6_ ( .D(n476), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[6]) );
  DFFRX1 MultResult_reg_reg_7_ ( .D(n477), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[7]) );
  DFFRX1 MultResult_reg_reg_8_ ( .D(n478), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[8]) );
  DFFRX1 MultResult_reg_reg_9_ ( .D(n479), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[9]) );
  DFFRX1 MultResult_reg_reg_10_ ( .D(n480), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[10]) );
  DFFRX1 MultResult_reg_reg_11_ ( .D(n481), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[11]) );
  DFFRX1 MultResult_reg_reg_12_ ( .D(n482), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[12]) );
  DFFRX1 MultResult_reg_reg_13_ ( .D(n483), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[13]) );
  DFFRX1 MultResult_reg_reg_14_ ( .D(n484), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[14]) );
  DFFRX1 MultResult_reg_reg_15_ ( .D(n485), .CLK(CLK), .CLRB(n408), .Q(
        MultResult_reg[15]) );
  DFFRX1 u_Adder_interconnect_Select_reg ( .D(n1723), .CLK(CLK), .CLRB(n408), 
        .Q(AddSelect) );
  FULLADD add_x_176_U9 ( .A(Add_Op1_wire[1]), .B(Add_Op2_wire[1]), .CIN(n1749), 
        .COUT(add_x_176_n12), .SUM(u_adder_24b_N123) );
  FULLADD add_x_176_U8 ( .A(Add_Op1_wire[2]), .B(Add_Op2_wire[2]), .CIN(
        add_x_176_n12), .COUT(add_x_176_n11), .SUM(u_adder_24b_N124) );
  FULLADD add_x_176_U7 ( .A(Add_Op1_wire[3]), .B(Add_Op2_wire[3]), .CIN(
        add_x_176_n11), .COUT(add_x_176_n10), .SUM(u_adder_24b_N125) );
  FULLADD add_x_176_U6 ( .A(Add_Op1_wire[4]), .B(Add_Op2_wire[4]), .CIN(
        add_x_176_n10), .COUT(add_x_176_n9), .SUM(u_adder_24b_N126) );
  FULLADD add_x_176_U5 ( .A(Add_Op1_wire[5]), .B(Add_Op2_wire[5]), .CIN(
        add_x_176_n9), .COUT(add_x_176_n8), .SUM(u_adder_24b_N127) );
  FULLADD add_x_176_U4 ( .A(Add_Op1_wire[6]), .B(Add_Op2_wire[6]), .CIN(
        add_x_176_n8), .COUT(add_x_176_n7), .SUM(u_adder_24b_N128) );
  FULLADD add_x_176_U3 ( .A(Add_Op1_wire[7]), .B(Add_Op2_wire[7]), .CIN(
        add_x_176_n7), .COUT(add_x_176_n6), .SUM(u_adder_24b_N129) );
  FULLADD add_x_176_U2 ( .A(Add_Op1_wire[8]), .B(Add_Op2_wire[8]), .CIN(n1750), 
        .COUT(u_adder_24b_N131), .SUM(u_adder_24b_N130) );
  BUF4X U1588 ( .IN(n1921), .OUT(n1819) );
  NAND3X1 U1589 ( .IN1(n1834), .IN2(Booth_valid), .IN3(n732), .OUT(n1725) );
  NAND2X1 U1590 ( .IN1(n1901), .IN2(n1725), .OUT(n1897) );
  INVX1 U1591 ( .IN(n1867), .OUT(n1726) );
  NOR2X1 U1592 ( .IN1(n2038), .IN2(n1726), .OUT(n1883) );
  NAND3X1 U1593 ( .IN1(n2053), .IN2(n1898), .IN3(Booth_Add_ack), .OUT(n1727)
         );
  INVX1 U1594 ( .IN(n1727), .OUT(n1903) );
  INVX1 U1595 ( .IN(n1890), .OUT(n1728) );
  NOR2X1 U1596 ( .IN1(Booth_valid), .IN2(n1728), .OUT(n1882) );
  AOI21 U1597 ( .IN1(n1898), .IN2(n1847), .IN3(n1889), .OUT(n1729) );
  NAND2X1 U1598 ( .IN1(n2104), .IN2(n1729), .OUT(n1556) );
  INVX4 U1599 ( .IN(AdderCntrl_ExcCheck_Datain[7]), .OUT(n1731) );
  INVX4 U1600 ( .IN(AdderCntrl_ExcCheck_Datain[10]), .OUT(n1732) );
  INVX4 U1601 ( .IN(n1834), .OUT(n1833) );
  INVX1 U1602 ( .IN(n2142), .OUT(n588) );
  INVX1 U1603 ( .IN(n2118), .OUT(n602) );
  INVX1 U1604 ( .IN(n2117), .OUT(n603) );
  INVX1 U1605 ( .IN(n2080), .OUT(n703) );
  INVX1 U1606 ( .IN(n2116), .OUT(n604) );
  INVX1 U1607 ( .IN(n2200), .OUT(n530) );
  INVX1 U1608 ( .IN(n2181), .OUT(n549) );
  INVX1 U1609 ( .IN(n2182), .OUT(n548) );
  INVX1 U1610 ( .IN(n2184), .OUT(n546) );
  INVX1 U1611 ( .IN(n2196), .OUT(n534) );
  INVX1 U1612 ( .IN(n2190), .OUT(n540) );
  INVX1 U1613 ( .IN(n2191), .OUT(n539) );
  INVX1 U1614 ( .IN(n2183), .OUT(n547) );
  INVX1 U1615 ( .IN(n2180), .OUT(n550) );
  INVX1 U1616 ( .IN(n2203), .OUT(n527) );
  INVX1 U1617 ( .IN(n2202), .OUT(n528) );
  INVX1 U1618 ( .IN(n2186), .OUT(n544) );
  INVX1 U1619 ( .IN(n2115), .OUT(n605) );
  INVX1 U1620 ( .IN(n2189), .OUT(n541) );
  INVX1 U1621 ( .IN(n2185), .OUT(n545) );
  INVX1 U1622 ( .IN(n2193), .OUT(n537) );
  INVX1 U1623 ( .IN(n2188), .OUT(n542) );
  INVX1 U1624 ( .IN(n2192), .OUT(n538) );
  INVX1 U1625 ( .IN(n2204), .OUT(n526) );
  INVX1 U1626 ( .IN(n2179), .OUT(n551) );
  INVX1 U1627 ( .IN(n2187), .OUT(n543) );
  INVX1 U1628 ( .IN(n2155), .OUT(n572) );
  INVX1 U1629 ( .IN(n2153), .OUT(n574) );
  INVX1 U1630 ( .IN(n2152), .OUT(n575) );
  INVX1 U1631 ( .IN(n2151), .OUT(n576) );
  INVX1 U1632 ( .IN(n2156), .OUT(n571) );
  INVX1 U1633 ( .IN(n2150), .OUT(n577) );
  INVX1 U1634 ( .IN(n2149), .OUT(n578) );
  INVX1 U1635 ( .IN(n2158), .OUT(n569) );
  INVX1 U1636 ( .IN(n2148), .OUT(n579) );
  INVX1 U1637 ( .IN(n2147), .OUT(n580) );
  INVX1 U1638 ( .IN(n2159), .OUT(n568) );
  INVX1 U1639 ( .IN(n2146), .OUT(n581) );
  INVX1 U1640 ( .IN(n2145), .OUT(n582) );
  INVX1 U1641 ( .IN(n2212), .OUT(n520) );
  INVX1 U1642 ( .IN(n2144), .OUT(n583) );
  INVX1 U1643 ( .IN(n2209), .OUT(n521) );
  INVX1 U1644 ( .IN(n2162), .OUT(n565) );
  INVX1 U1645 ( .IN(n2208), .OUT(n522) );
  INVX1 U1646 ( .IN(n2163), .OUT(n564) );
  INVX1 U1647 ( .IN(n2164), .OUT(n563) );
  INVX1 U1648 ( .IN(n2154), .OUT(n573) );
  INVX1 U1649 ( .IN(n2207), .OUT(n523) );
  INVX1 U1650 ( .IN(n2171), .OUT(n556) );
  INVX1 U1651 ( .IN(n2177), .OUT(n552) );
  INVX1 U1652 ( .IN(n2170), .OUT(n557) );
  INVX1 U1653 ( .IN(n2167), .OUT(n560) );
  INVX1 U1654 ( .IN(n2172), .OUT(n555) );
  INVX1 U1655 ( .IN(n2168), .OUT(n559) );
  INVX1 U1656 ( .IN(n2205), .OUT(n525) );
  INVX1 U1657 ( .IN(n2206), .OUT(n524) );
  INVX1 U1658 ( .IN(n2169), .OUT(n558) );
  INVX1 U1659 ( .IN(n2173), .OUT(n554) );
  INVX1 U1660 ( .IN(n2084), .OUT(n702) );
  INVX1 U1661 ( .IN(n2088), .OUT(n701) );
  INVX1 U1662 ( .IN(n2092), .OUT(n700) );
  INVX1 U1663 ( .IN(n2096), .OUT(n699) );
  INVX1 U1664 ( .IN(n2174), .OUT(n553) );
  INVX1 U1665 ( .IN(n2077), .OUT(n2078) );
  INVX1 U1666 ( .IN(n2166), .OUT(n561) );
  INVX1 U1667 ( .IN(n2165), .OUT(n562) );
  INVX1 U1668 ( .IN(n2161), .OUT(n566) );
  INVX1 U1669 ( .IN(n2160), .OUT(n567) );
  INVX1 U1670 ( .IN(n2157), .OUT(n570) );
  INVX1 U1671 ( .IN(n2198), .OUT(n532) );
  INVX1 U1672 ( .IN(n2194), .OUT(n536) );
  INVX1 U1673 ( .IN(n2199), .OUT(n531) );
  INVX1 U1674 ( .IN(n2201), .OUT(n529) );
  INVX1 U1675 ( .IN(n2125), .OUT(n596) );
  INVX1 U1676 ( .IN(n2197), .OUT(n533) );
  INVX1 U1677 ( .IN(n2195), .OUT(n535) );
  INVX1 U1678 ( .IN(n2242), .OUT(n426) );
  INVX1 U1679 ( .IN(n2245), .OUT(n423) );
  INVX1 U1680 ( .IN(n2255), .OUT(n413) );
  INVX1 U1681 ( .IN(n2254), .OUT(n414) );
  INVX1 U1682 ( .IN(n2243), .OUT(n425) );
  INVX1 U1683 ( .IN(n2244), .OUT(n424) );
  INVX1 U1684 ( .IN(n2241), .OUT(n427) );
  INVX1 U1685 ( .IN(n2258), .OUT(n412) );
  INVX1 U1686 ( .IN(n2246), .OUT(n422) );
  INVX1 U1687 ( .IN(n2253), .OUT(n415) );
  INVX1 U1688 ( .IN(n2240), .OUT(n428) );
  INVX1 U1689 ( .IN(n2252), .OUT(n416) );
  INVX4 U1690 ( .IN(n2211), .OUT(n1832) );
  INVX1 U1691 ( .IN(n2251), .OUT(n417) );
  INVX1 U1692 ( .IN(n2247), .OUT(n421) );
  INVX1 U1693 ( .IN(n2250), .OUT(n418) );
  INVX1 U1694 ( .IN(n2249), .OUT(n419) );
  NANDX2 U1695 ( .IN1(n1796), .IN2(n1895), .OUT(n2056) );
  INVX1 U1696 ( .IN(n2248), .OUT(n420) );
  INVX1 U1697 ( .IN(n2221), .OUT(n479) );
  INVX1 U1698 ( .IN(n2235), .OUT(n467) );
  INVX1 U1699 ( .IN(n2220), .OUT(n480) );
  INVX1 U1700 ( .IN(n2232), .OUT(n468) );
  INVX1 U1701 ( .IN(n2222), .OUT(n478) );
  INVX1 U1702 ( .IN(n2231), .OUT(n469) );
  INVX1 U1703 ( .IN(n2230), .OUT(n470) );
  INVX1 U1704 ( .IN(n2219), .OUT(n481) );
  INVX1 U1705 ( .IN(n2218), .OUT(n482) );
  INVX1 U1706 ( .IN(n2229), .OUT(n471) );
  INVX1 U1707 ( .IN(n2217), .OUT(n483) );
  INVX1 U1708 ( .IN(n2216), .OUT(n484) );
  NAND2X1 U1709 ( .IN1(n2016), .IN2(n2015), .OUT(n2017) );
  INVX1 U1710 ( .IN(n2223), .OUT(n477) );
  INVX1 U1711 ( .IN(n2215), .OUT(n485) );
  INVX1 U1712 ( .IN(n2224), .OUT(n476) );
  INVX1 U1713 ( .IN(n2226), .OUT(n474) );
  INVX1 U1714 ( .IN(n2228), .OUT(n472) );
  INVX1 U1715 ( .IN(n2225), .OUT(n475) );
  INVX4 U1716 ( .IN(n2175), .OUT(n1826) );
  INVX1 U1717 ( .IN(n2227), .OUT(n473) );
  NANDX2 U1718 ( .IN1(n1800), .IN2(n1862), .OUT(n1850) );
  INVX1 U1719 ( .IN(n2111), .OUT(n611) );
  NANDX2 U1720 ( .IN1(n1801), .IN2(n1862), .OUT(n1863) );
  INVX1 U1721 ( .IN(n2114), .OUT(n610) );
  NAND2X1 U1722 ( .IN1(n1840), .IN2(n1896), .OUT(n1839) );
  NAND2X1 U1723 ( .IN1(n2011), .IN2(n2010), .OUT(n2012) );
  INVX1 U1724 ( .IN(n2081), .OUT(n2082) );
  NANDX2 U1725 ( .IN1(n1797), .IN2(n1862), .OUT(n1853) );
  NANDX2 U1726 ( .IN1(n1799), .IN2(n1862), .OUT(n1859) );
  NANDX2 U1727 ( .IN1(n1798), .IN2(n1862), .OUT(n1856) );
  INVX1 U1728 ( .IN(n2105), .OUT(n617) );
  NANDX2 U1729 ( .IN1(Booth_Add_datain1[8]), .IN2(n1803), .OUT(n1913) );
  INVX1 U1730 ( .IN(n2106), .OUT(n616) );
  INVX1 U1731 ( .IN(MulCntrl_ExcCheck_Datain[13]), .OUT(n2002) );
  INVX1 U1732 ( .IN(n2110), .OUT(n612) );
  INVX1 U1733 ( .IN(n2109), .OUT(n613) );
  NAND2X1 U1734 ( .IN1(n1894), .IN2(n2101), .OUT(n1895) );
  INVX1 U1735 ( .IN(n2108), .OUT(n614) );
  NAND2X1 U1736 ( .IN1(MulCntrl_ExcCheck_Datain[12]), .IN2(
        MulCntrl_ExcCheck_Datain[11]), .OUT(n2000) );
  INVX1 U1737 ( .IN(n2107), .OUT(n615) );
  INVX1 U1738 ( .IN(n1940), .OUT(DEBUG[4]) );
  INVX1 U1739 ( .IN(n1937), .OUT(DEBUG[3]) );
  INVX1 U1740 ( .IN(n1936), .OUT(DEBUG[2]) );
  INVX1 U1741 ( .IN(Add_Op1_wire[0]), .OUT(n1747) );
  NAND2X1 U1742 ( .IN1(n2236), .IN2(n2213), .OUT(N193) );
  INVX1 U1743 ( .IN(n1897), .OUT(n1894) );
  INVX1 U1744 ( .IN(n2239), .OUT(n429) );
  INVX1 U1745 ( .IN(n2238), .OUT(n430) );
  INVX4 U1746 ( .IN(n1816), .OUT(Booth_ack) );
  INVX1 U1747 ( .IN(n1950), .OUT(DOUT[2]) );
  INVX1 U1748 ( .IN(n1948), .OUT(DOUT[15]) );
  INVX1 U1749 ( .IN(n1944), .OUT(DOUT[11]) );
  INVX1 U1750 ( .IN(n1957), .OUT(DOUT[9]) );
  INVX1 U1751 ( .IN(n1946), .OUT(DOUT[13]) );
  INVX1 U1752 ( .IN(n1949), .OUT(DOUT[1]) );
  INVX1 U1753 ( .IN(n1947), .OUT(DOUT[14]) );
  INVX1 U1754 ( .IN(n1958), .OUT(DOV) );
  INVX1 U1755 ( .IN(AdderCntrl_ExcCheck_Datain[13]), .OUT(n2020) );
  INVX1 U1756 ( .IN(n1945), .OUT(DOUT[12]) );
  INVX1 U1757 ( .IN(n1942), .OUT(DOUT[0]) );
  INVX1 U1758 ( .IN(n1956), .OUT(DOUT[8]) );
  NANDX2 U1759 ( .IN1(n1779), .IN2(n1885), .OUT(n1835) );
  INVX1 U1760 ( .IN(n1953), .OUT(DOUT[5]) );
  INVX1 U1761 ( .IN(n1954), .OUT(DOUT[6]) );
  INVX1 U1762 ( .IN(n1959), .OUT(EXC[0]) );
  INVX1 U1763 ( .IN(n1952), .OUT(DOUT[4]) );
  INVX1 U1764 ( .IN(n1960), .OUT(EXC[1]) );
  INVX1 U1765 ( .IN(n1955), .OUT(DOUT[7]) );
  INVX4 U1766 ( .IN(n2210), .OUT(n1830) );
  INVX1 U1767 ( .IN(n1961), .OUT(EXC[2]) );
  INVX1 U1768 ( .IN(n2085), .OUT(n2086) );
  INVX4 U1769 ( .IN(n2176), .OUT(n1828) );
  INVX1 U1770 ( .IN(n1951), .OUT(DOUT[3]) );
  NANDX2 U1771 ( .IN1(n1766), .IN2(n1898), .OUT(n1899) );
  INVX1 U1772 ( .IN(n1928), .OUT(DACK) );
  INVX1 U1773 ( .IN(n1943), .OUT(DOUT[10]) );
  INVX1 U1774 ( .IN(n1997), .OUT(n1656) );
  INVX1 U1775 ( .IN(n2052), .OUT(n1587) );
  INVX1 U1776 ( .IN(n2130), .OUT(n594) );
  INVX1 U1777 ( .IN(n2135), .OUT(n592) );
  INVX1 U1778 ( .IN(n1847), .OUT(n1848) );
  INVX1 U1779 ( .IN(n2139), .OUT(n2140) );
  INVX1 U1780 ( .IN(u_exc_check_N45), .OUT(n2102) );
  INVX1 U1781 ( .IN(n2089), .OUT(n2090) );
  INVX1 U1782 ( .IN(n2094), .OUT(n2093) );
  INVX1 U1783 ( .IN(n2131), .OUT(n2133) );
  INVX1 U1784 ( .IN(n2126), .OUT(n2129) );
  INVX1 U1785 ( .IN(n2068), .OUT(n1996) );
  INVX1 U1786 ( .IN(n2066), .OUT(n2051) );
  BUF4X U1787 ( .IN(AdderCntrl_Op1[7]), .OUT(n1808) );
  NANDX2 U1788 ( .IN1(n462), .IN2(n1764), .OUT(n1975) );
  NANDX2 U1789 ( .IN1(n1834), .IN2(u_booth_BStateMC_1_), .OUT(n1901) );
  NANDX2 U1790 ( .IN1(multStateMC[0]), .IN2(n1755), .OUT(n1976) );
  INVX1 U1791 ( .IN(n1929), .OUT(n1935) );
  INVX4 U1792 ( .IN(CS), .OUT(n2061) );
  INVX4 U1793 ( .IN(n1736), .OUT(n1739) );
  INVX4 U1794 ( .IN(n1733), .OUT(n1740) );
  INVX4 U1795 ( .IN(n1741), .OUT(n1742) );
  INVX4 U1796 ( .IN(n1743), .OUT(n1744) );
  INVX4 U1797 ( .IN(n1745), .OUT(n1746) );
  MUX2X1 U1798 ( .IN1(n1747), .IN2(Add_Op1_wire[0]), .S(n1748), .OUT(
        u_adder_24b_N122) );
  NOR2X1 U1799 ( .IN1(n1747), .IN2(n1748), .OUT(add_x_176_n13) );
  BUF4X U1800 ( .IN(add_x_176_n13), .OUT(n1749) );
  BUF4X U1801 ( .IN(add_x_176_n6), .OUT(n1750) );
  INVX4 U1802 ( .IN(Add_Op2_wire[0]), .OUT(n1748) );
  INVX1 U1803 ( .IN(n2123), .OUT(n597) );
  BUF4X U1804 ( .IN(n1888), .OUT(n1816) );
  INVX4 U1805 ( .IN(n1826), .OUT(n1825) );
  INVX4 U1806 ( .IN(n1832), .OUT(n1831) );
  INVX4 U1807 ( .IN(n1830), .OUT(n1829) );
  NANDX2 U1808 ( .IN1(n695), .IN2(n694), .OUT(n1846) );
  BUF4X U1809 ( .IN(AdderCntrl_Op2[8]), .OUT(n1809) );
  NANDX2 U1810 ( .IN1(n1905), .IN2(n1898), .OUT(n1849) );
  BUF4X U1811 ( .IN(n1819), .OUT(n1802) );
  NANDX2 U1812 ( .IN1(n1902), .IN2(n2058), .OUT(n1546) );
  NANDX2 U1813 ( .IN1(n1852), .IN2(n1851), .OUT(n1549) );
  NANDX2 U1814 ( .IN1(n1855), .IN2(n1854), .OUT(n1550) );
  NAND2X1 U1815 ( .IN1(n1834), .IN2(n1867), .OUT(n1836) );
  NANDX2 U1816 ( .IN1(n2057), .IN2(n2056), .OUT(n1547) );
  NANDX2 U1817 ( .IN1(n2055), .IN2(n2054), .OUT(n1548) );
  NANDX2 U1818 ( .IN1(n1865), .IN2(n1864), .OUT(n1553) );
  NANDX2 U1819 ( .IN1(n1861), .IN2(n1860), .OUT(n1552) );
  NANDX2 U1820 ( .IN1(n1858), .IN2(n1857), .OUT(n1551) );
  NANDX2 U1821 ( .IN1(n1834), .IN2(n2059), .OUT(n2060) );
  NANDX2 U1822 ( .IN1(n1834), .IN2(n2064), .OUT(n992) );
  BUF4X U1823 ( .IN(n2256), .OUT(n1824) );
  BUF4X U1824 ( .IN(n2233), .OUT(n1823) );
  BUF4X U1825 ( .IN(n1971), .OUT(n1821) );
  BUF4X U1826 ( .IN(n1974), .OUT(n1820) );
  NANDX2 U1827 ( .IN1(u_exc_check_N45), .IN2(n2036), .OUT(n2037) );
  BUF4X U1828 ( .IN(n2124), .OUT(n1822) );
  INVX1 U1829 ( .IN(MODE[2]), .OUT(n1932) );
  NANDX2 U1830 ( .IN1(n1834), .IN2(n1982), .OUT(n1302) );
  NANDX2 U1831 ( .IN1(n1834), .IN2(n1882), .OUT(n2104) );
  INVX4 U1832 ( .IN(n1850), .OUT(u_booth_N53) );
  INVX4 U1833 ( .IN(n1853), .OUT(u_booth_N52) );
  INVX4 U1834 ( .IN(n1863), .OUT(u_booth_N49) );
  INVX4 U1835 ( .IN(n1859), .OUT(u_booth_N50) );
  INVX4 U1836 ( .IN(n1856), .OUT(u_booth_N51) );
  INVX4 U1837 ( .IN(n1843), .OUT(n1893) );
  NAND2X1 U1838 ( .IN1(RSTn), .IN2(n1972), .OUT(n1973) );
  NAND2X1 U1839 ( .IN1(n587), .IN2(CS), .OUT(n1941) );
  INVX4 U1840 ( .IN(n2075), .OUT(n2097) );
  INVX4 U1841 ( .IN(n2053), .OUT(n1905) );
  NANDX2 U1842 ( .IN1(n1837), .IN2(n1898), .OUT(n1843) );
  NANDX2 U1843 ( .IN1(n2072), .IN2(n2071), .OUT(n2076) );
  INVX4 U1844 ( .IN(n1899), .OUT(n2072) );
  INVX4 U1845 ( .IN(n2137), .OUT(n2035) );
  NANDX2 U1846 ( .IN1(n2025), .IN2(n2030), .OUT(n2137) );
  NANDX2 U1847 ( .IN1(RSTn), .IN2(n1998), .OUT(n2139) );
  INVX4 U1848 ( .IN(n1914), .OUT(Add_Op2_wire[1]) );
  INVX4 U1849 ( .IN(n1906), .OUT(Add_Op1_wire[1]) );
  INVX4 U1850 ( .IN(n1915), .OUT(Add_Op2_wire[2]) );
  INVX4 U1851 ( .IN(n1907), .OUT(Add_Op1_wire[2]) );
  INVX4 U1852 ( .IN(n1916), .OUT(Add_Op2_wire[3]) );
  INVX4 U1853 ( .IN(n1908), .OUT(Add_Op1_wire[3]) );
  INVX4 U1854 ( .IN(n1917), .OUT(Add_Op2_wire[4]) );
  INVX4 U1855 ( .IN(n1909), .OUT(Add_Op1_wire[4]) );
  INVX4 U1856 ( .IN(n1918), .OUT(Add_Op2_wire[5]) );
  INVX4 U1857 ( .IN(n1910), .OUT(Add_Op1_wire[5]) );
  INVX4 U1858 ( .IN(n1919), .OUT(Add_Op2_wire[6]) );
  INVX4 U1859 ( .IN(n1911), .OUT(Add_Op1_wire[6]) );
  INVX4 U1860 ( .IN(n1920), .OUT(Add_Op2_wire[7]) );
  INVX4 U1861 ( .IN(n1912), .OUT(Add_Op1_wire[7]) );
  INVX4 U1862 ( .IN(n1922), .OUT(Add_Op2_wire[8]) );
  INVX4 U1863 ( .IN(n1913), .OUT(Add_Op1_wire[8]) );
  INVX4 U1864 ( .IN(n1806), .OUT(n1803) );
  NANDX2 U1865 ( .IN1(n1759), .IN2(n1807), .OUT(n1806) );
  INVX4 U1866 ( .IN(n1819), .OUT(n1807) );
  INVX4 U1867 ( .IN(n1811), .OUT(n1812) );
  INVX4 U1868 ( .IN(n1752), .OUT(n1815) );
  BUF4X U1869 ( .IN(AdderCntrl_Op1[8]), .OUT(n1810) );
  BUF4X U1870 ( .IN(RSTn), .OUT(n1834) );
  NAND2X1 U1871 ( .IN1(RSTn), .IN2(n1969), .OUT(n1970) );
  NAND2X1 U1872 ( .IN1(u_booth_count_reg_2_), .IN2(n1892), .OUT(n1841) );
  BUF4X U1873 ( .IN(MulCntrl_Op1[13]), .OUT(n1814) );
  NAND2X1 U1874 ( .IN1(n1795), .IN2(n1895), .OUT(n2054) );
  INVX4 U1875 ( .IN(n2104), .OUT(n2112) );
  INVX4 U1876 ( .IN(n2076), .OUT(n2098) );
  NAND2X1 U1877 ( .IN1(n1834), .IN2(n1835), .OUT(n1896) );
  NAND2X1 U1878 ( .IN1(n2053), .IN2(n1766), .OUT(n1837) );
  INVX4 U1879 ( .IN(n1975), .OUT(n2237) );
  INVX4 U1880 ( .IN(n1976), .OUT(n2214) );
  NAND2X1 U1881 ( .IN1(Add_Op2[0]), .IN2(n1819), .OUT(n1804) );
  NAND2X1 U1882 ( .IN1(Add_Op1[0]), .IN2(n1819), .OUT(n1805) );
  INVX4 U1883 ( .IN(n1751), .OUT(n1818) );
  INVX4 U1884 ( .IN(n1813), .OUT(n1817) );
  INVX4 U1885 ( .IN(n1828), .OUT(n1827) );
  AOI22 U1886 ( .IN1(Add_Op2[1]), .IN2(n1819), .IN3(Booth_Add_datain2[1]), 
        .IN4(n1803), .OUT(n1914) );
  AOI22 U1887 ( .IN1(Add_Op1[1]), .IN2(n1819), .IN3(Booth_Add_datain1[1]), 
        .IN4(n1803), .OUT(n1906) );
  AOI22 U1888 ( .IN1(Add_Op2[2]), .IN2(n1802), .IN3(Booth_Add_datain2[2]), 
        .IN4(n1803), .OUT(n1915) );
  AOI22 U1889 ( .IN1(Add_Op1[2]), .IN2(n1802), .IN3(Booth_Add_datain1[2]), 
        .IN4(n1803), .OUT(n1907) );
  AOI22 U1890 ( .IN1(Add_Op2[3]), .IN2(n1802), .IN3(Booth_Add_datain2[3]), 
        .IN4(n1803), .OUT(n1916) );
  AOI22 U1891 ( .IN1(Add_Op1[3]), .IN2(n1802), .IN3(Booth_Add_datain1[3]), 
        .IN4(n1803), .OUT(n1908) );
  AOI22 U1892 ( .IN1(Add_Op2[4]), .IN2(n1802), .IN3(Booth_Add_datain2[4]), 
        .IN4(n1803), .OUT(n1917) );
  AOI22 U1893 ( .IN1(Add_Op1[4]), .IN2(n1802), .IN3(Booth_Add_datain1[4]), 
        .IN4(n1803), .OUT(n1909) );
  AOI22 U1894 ( .IN1(Add_Op2[5]), .IN2(n1802), .IN3(Booth_Add_datain2[5]), 
        .IN4(n1803), .OUT(n1918) );
  AOI22 U1895 ( .IN1(Add_Op1[5]), .IN2(n1802), .IN3(Booth_Add_datain1[5]), 
        .IN4(n1803), .OUT(n1910) );
  AOI22 U1896 ( .IN1(Add_Op2[6]), .IN2(n1802), .IN3(Booth_Add_datain2[6]), 
        .IN4(n1803), .OUT(n1919) );
  AOI22 U1897 ( .IN1(Add_Op1[6]), .IN2(n1802), .IN3(Booth_Add_datain1[6]), 
        .IN4(n1803), .OUT(n1911) );
  AOI22 U1898 ( .IN1(Add_Op2[7]), .IN2(n1802), .IN3(Booth_Add_datain2[7]), 
        .IN4(n1803), .OUT(n1920) );
  AOI22 U1899 ( .IN1(Add_Op1[7]), .IN2(n1802), .IN3(Booth_Add_datain1[7]), 
        .IN4(n1803), .OUT(n1912) );
  AOI22 U1900 ( .IN1(Add_Op2[8]), .IN2(n1802), .IN3(Booth_Add_datain2[8]), 
        .IN4(n1803), .OUT(n1922) );
  OAI21 U1901 ( .IN1(n1760), .IN2(n1806), .IN3(n1804), .OUT(Add_Op2_wire[0])
         );
  OAI21 U1902 ( .IN1(n1758), .IN2(n1806), .IN3(n1805), .OUT(Add_Op1_wire[0])
         );
  TIEHI U1903 ( .OUT(n408) );
  NAND2X1 U1904 ( .IN1(u_booth_count_reg_2_), .IN2(n1840), .OUT(n1844) );
  INVX4 U1905 ( .IN(n2070), .OUT(u_adder_24b_N52) );
  INVX4 U1906 ( .IN(n2213), .OUT(n2234) );
  INVX4 U1907 ( .IN(n2236), .OUT(n2257) );
  NOR2X1 U1908 ( .IN1(n732), .IN2(u_booth_BStateMC_1_), .OUT(n1867) );
  NOR2X1 U1909 ( .IN1(u_booth_BStateMC_1_), .IN2(n1765), .OUT(n1890) );
  AOI22 U1910 ( .IN1(n1867), .IN2(n2038), .IN3(Booth_valid), .IN4(n1890), 
        .OUT(n1885) );
  INVX4 U1911 ( .IN(n1896), .OUT(n1892) );
  INVX4 U1912 ( .IN(n1836), .OUT(n1898) );
  MUX2X1 U1913 ( .IN1(n1892), .IN2(n1893), .S(n694), .OUT(n1554) );
  NOR2X1 U1914 ( .IN1(n694), .IN2(n695), .OUT(n1840) );
  OAI21 U1915 ( .IN1(n695), .IN2(n1896), .IN3(n1843), .OUT(n1838) );
  NAND3X1 U1916 ( .IN1(n1846), .IN2(n1839), .IN3(n1838), .OUT(n1079) );
  OAI21 U1917 ( .IN1(n1840), .IN2(u_booth_count_reg_2_), .IN3(n1844), .OUT(
        n1842) );
  OAI21 U1918 ( .IN1(n1843), .IN2(n1842), .IN3(n1841), .OUT(n1555) );
  MUX2X1 U1919 ( .IN1(n1789), .IN2(u_booth_count_reg_3_), .S(n1844), .OUT(
        n1845) );
  AOI22 U1920 ( .IN1(n1893), .IN2(n1845), .IN3(u_booth_count_reg_3_), .IN4(
        n1892), .OUT(n1092) );
  NOR2X1 U1921 ( .IN1(n732), .IN2(n1901), .OUT(n1889) );
  OAI21 U1922 ( .IN1(u_booth_count_reg_2_), .IN2(n1846), .IN3(
        u_booth_count_reg_3_), .OUT(n1847) );
  NANDX2 U1923 ( .IN1(n1867), .IN2(n1848), .OUT(n1888) );
  AOI21 U1924 ( .IN1(Booth_ack), .IN2(n1834), .IN3(n1889), .OUT(n1088) );
  NANDX2 U1925 ( .IN1(n2038), .IN2(n1898), .OUT(n2101) );
  AOI22 U1926 ( .IN1(n1800), .IN2(n1897), .IN3(Add_dataout[5]), .IN4(n1903), 
        .OUT(n1852) );
  INVX4 U1927 ( .IN(n1849), .OUT(n1904) );
  INVX4 U1928 ( .IN(n2101), .OUT(n1862) );
  AOI21 U1929 ( .IN1(n1904), .IN2(n1795), .IN3(u_booth_N53), .OUT(n1851) );
  AOI22 U1930 ( .IN1(n1897), .IN2(n1797), .IN3(Add_dataout[4]), .IN4(n1903), 
        .OUT(n1855) );
  AOI21 U1931 ( .IN1(n1904), .IN2(n1800), .IN3(u_booth_N52), .OUT(n1854) );
  AOI22 U1932 ( .IN1(n1897), .IN2(n1798), .IN3(Add_dataout[3]), .IN4(n1903), 
        .OUT(n1858) );
  AOI21 U1933 ( .IN1(n1904), .IN2(n1797), .IN3(u_booth_N51), .OUT(n1857) );
  AOI22 U1934 ( .IN1(n1897), .IN2(n1799), .IN3(Add_dataout[2]), .IN4(n1903), 
        .OUT(n1861) );
  AOI21 U1935 ( .IN1(n1904), .IN2(n1798), .IN3(u_booth_N50), .OUT(n1860) );
  AOI22 U1936 ( .IN1(n1801), .IN2(n1897), .IN3(Add_dataout[1]), .IN4(n1903), 
        .OUT(n1865) );
  AOI21 U1937 ( .IN1(n1904), .IN2(n1799), .IN3(u_booth_N49), .OUT(n1864) );
  AOI22 U1938 ( .IN1(n1904), .IN2(n1801), .IN3(n1903), .IN4(Add_dataout[0]), 
        .OUT(n1866) );
  OAI21 U1939 ( .IN1(n721), .IN2(n1896), .IN3(n1866), .OUT(n1544) );
  INVX4 U1940 ( .IN(n1901), .OUT(n1887) );
  AOI22 U1941 ( .IN1(n1883), .IN2(n1790), .IN3(Booth_datain2[7]), .IN4(n1882), 
        .OUT(n1868) );
  OAI21 U1942 ( .IN1(n1885), .IN2(n720), .IN3(n1868), .OUT(n1869) );
  AOI22 U1943 ( .IN1(n1887), .IN2(n1781), .IN3(n1834), .IN4(n1869), .OUT(n1022) );
  AOI22 U1944 ( .IN1(n1883), .IN2(n1781), .IN3(Booth_datain2[6]), .IN4(n1882), 
        .OUT(n1870) );
  OAI21 U1945 ( .IN1(n1885), .IN2(n719), .IN3(n1870), .OUT(n1871) );
  AOI22 U1946 ( .IN1(n1887), .IN2(n1782), .IN3(n1834), .IN4(n1871), .OUT(n1028) );
  AOI22 U1947 ( .IN1(n1883), .IN2(n1782), .IN3(Booth_datain2[5]), .IN4(n1882), 
        .OUT(n1872) );
  OAI21 U1948 ( .IN1(n1885), .IN2(n718), .IN3(n1872), .OUT(n1873) );
  AOI22 U1949 ( .IN1(n1887), .IN2(n1783), .IN3(RSTn), .IN4(n1873), .OUT(n1031)
         );
  AOI22 U1950 ( .IN1(n1883), .IN2(n1783), .IN3(Booth_datain2[4]), .IN4(n1882), 
        .OUT(n1874) );
  OAI21 U1951 ( .IN1(n1885), .IN2(n717), .IN3(n1874), .OUT(n1875) );
  AOI22 U1952 ( .IN1(n1887), .IN2(n1784), .IN3(RSTn), .IN4(n1875), .OUT(n1034)
         );
  AOI22 U1953 ( .IN1(n1883), .IN2(n1784), .IN3(Booth_datain2[3]), .IN4(n1882), 
        .OUT(n1876) );
  OAI21 U1954 ( .IN1(n1885), .IN2(n716), .IN3(n1876), .OUT(n1877) );
  AOI22 U1955 ( .IN1(n1887), .IN2(n1785), .IN3(RSTn), .IN4(n1877), .OUT(n1037)
         );
  AOI22 U1956 ( .IN1(n1883), .IN2(n1785), .IN3(Booth_datain2[2]), .IN4(n1882), 
        .OUT(n1878) );
  OAI21 U1957 ( .IN1(n1885), .IN2(n715), .IN3(n1878), .OUT(n1879) );
  AOI22 U1958 ( .IN1(n1887), .IN2(n1786), .IN3(RSTn), .IN4(n1879), .OUT(n1040)
         );
  AOI22 U1959 ( .IN1(n1883), .IN2(n1786), .IN3(Booth_datain2[1]), .IN4(n1882), 
        .OUT(n1880) );
  OAI21 U1960 ( .IN1(n1885), .IN2(n714), .IN3(n1880), .OUT(n1881) );
  AOI22 U1961 ( .IN1(n1887), .IN2(n1787), .IN3(RSTn), .IN4(n1881), .OUT(n1043)
         );
  AOI22 U1962 ( .IN1(n1883), .IN2(n1787), .IN3(Booth_datain2[0]), .IN4(n1882), 
        .OUT(n1884) );
  OAI21 U1963 ( .IN1(n1885), .IN2(n713), .IN3(n1884), .OUT(n1886) );
  AOI22 U1964 ( .IN1(n1887), .IN2(n1753), .IN3(RSTn), .IN4(n1886), .OUT(n1135)
         );
  NOR2X1 U1965 ( .IN1(n713), .IN2(n1816), .OUT(Booth_dataout[0]) );
  NOR2X1 U1966 ( .IN1(n714), .IN2(n1816), .OUT(Booth_dataout[1]) );
  NOR2X1 U1967 ( .IN1(n715), .IN2(n1816), .OUT(Booth_dataout[2]) );
  NOR2X1 U1968 ( .IN1(n716), .IN2(n1816), .OUT(Booth_dataout[3]) );
  NOR2X1 U1969 ( .IN1(n717), .IN2(n1816), .OUT(Booth_dataout[4]) );
  NOR2X1 U1970 ( .IN1(n718), .IN2(n1816), .OUT(Booth_dataout[5]) );
  NOR2X1 U1971 ( .IN1(n719), .IN2(n1816), .OUT(Booth_dataout[6]) );
  NOR2X1 U1972 ( .IN1(n720), .IN2(n1888), .OUT(Booth_dataout[7]) );
  NOR2X1 U1973 ( .IN1(n721), .IN2(n1888), .OUT(Booth_dataout[8]) );
  NOR2X1 U1974 ( .IN1(n722), .IN2(n1888), .OUT(Booth_dataout[9]) );
  NOR2X1 U1975 ( .IN1(n723), .IN2(n1888), .OUT(Booth_dataout[10]) );
  NOR2X1 U1976 ( .IN1(n724), .IN2(n1888), .OUT(Booth_dataout[11]) );
  NOR2X1 U1977 ( .IN1(n725), .IN2(n1888), .OUT(Booth_dataout[12]) );
  NOR2X1 U1978 ( .IN1(n726), .IN2(n1888), .OUT(Booth_dataout[13]) );
  NOR2X1 U1979 ( .IN1(n727), .IN2(n1816), .OUT(Booth_dataout[14]) );
  NOR2X1 U1980 ( .IN1(n728), .IN2(n1816), .OUT(Booth_dataout[15]) );
  AOI21 U1981 ( .IN1(n1890), .IN2(n1834), .IN3(n1889), .OUT(n1891) );
  OAI21 U1982 ( .IN1(n1891), .IN2(n1780), .IN3(n2101), .OUT(n1653) );
  AOI22 U1983 ( .IN1(n1893), .IN2(n1753), .IN3(u_booth_Q1_reg), .IN4(n1892), 
        .OUT(n1077) );
  AOI22 U1984 ( .IN1(n1904), .IN2(u_booth_A_reg_8_), .IN3(n1903), .IN4(
        Add_dataout[8]), .OUT(n1902) );
  OAI21 U1985 ( .IN1(n1896), .IN2(n1793), .IN3(n1902), .OUT(n1545) );
  NOR2X1 U1986 ( .IN1(n1776), .IN2(n2101), .OUT(n706) );
  AOI21 U1987 ( .IN1(u_booth_A_reg_7_), .IN2(n1897), .IN3(n706), .OUT(n2058)
         );
  OAI21 U1988 ( .IN1(Booth_valid), .IN2(n1765), .IN3(n1834), .OUT(n1900) );
  NANDX2 U1989 ( .IN1(n1901), .IN2(n1900), .OUT(n2113) );
  NOR2X1 U1990 ( .IN1(n728), .IN2(n2101), .OUT(u_booth_N55) );
  NOR2X1 U1991 ( .IN1(n727), .IN2(n2101), .OUT(u_booth_N54) );
  NOR2X1 U1992 ( .IN1(AddSelect), .IN2(n802), .OUT(n1921) );
  NAND3X1 U1993 ( .IN1(getdataStat_reg[0]), .IN2(n463), .IN3(ABUSY), .OUT(
        n1923) );
  NOR2X1 U1994 ( .IN1(n1923), .IN2(n1761), .OUT(AdderCntrl_valid) );
  NOR2X1 U1995 ( .IN1(ABUSY), .IN2(OPT), .OUT(n1924) );
  NAND3X1 U1996 ( .IN1(CS), .IN2(DIV), .IN3(n1924), .OUT(n1925) );
  NOR2X1 U1997 ( .IN1(getdataStat_reg[0]), .IN2(n1925), .OUT(n2178) );
  NOR2X1 U1998 ( .IN1(MBUSY), .IN2(getdataStat_reg[1]), .OUT(n1926) );
  NAND3X1 U1999 ( .IN1(DIV), .IN2(OPT), .IN3(n1926), .OUT(n1927) );
  NOR2X1 U2000 ( .IN1(n2061), .IN2(n1927), .OUT(n2143) );
  NOR2X1 U2001 ( .IN1(n2178), .IN2(n2143), .OUT(n1928) );
  NOR2X1 U2002 ( .IN1(MODE[1]), .IN2(MODE[0]), .OUT(n1929) );
  AOI22 U2003 ( .IN1(MODE[2]), .IN2(multStateMC[0]), .IN3(n1764), .IN4(n1932), 
        .OUT(n1931) );
  NOR2X1 U2004 ( .IN1(n1929), .IN2(MODE[2]), .OUT(n1939) );
  NOR2X1 U2005 ( .IN1(n1929), .IN2(n1932), .OUT(n1938) );
  AOI22 U2006 ( .IN1(n1939), .IN2(AdderCntrl_Debug[0]), .IN3(n1938), .IN4(
        MulCntrl_Debug[0]), .OUT(n1930) );
  OAI21 U2007 ( .IN1(n1935), .IN2(n1931), .IN3(n1930), .OUT(DEBUG[0]) );
  AOI22 U2008 ( .IN1(MODE[2]), .IN2(multStateMC[1]), .IN3(n1761), .IN4(n1932), 
        .OUT(n1934) );
  AOI22 U2009 ( .IN1(n1939), .IN2(AdderCntrl_Debug[1]), .IN3(n1938), .IN4(
        MulCntrl_Debug[1]), .OUT(n1933) );
  OAI21 U2010 ( .IN1(n1935), .IN2(n1934), .IN3(n1933), .OUT(DEBUG[1]) );
  AOI22 U2011 ( .IN1(n1939), .IN2(AdderCntrl_Debug[2]), .IN3(n1938), .IN4(
        MulCntrl_Debug[2]), .OUT(n1936) );
  AOI22 U2012 ( .IN1(n1939), .IN2(AdderCntrl_Debug[3]), .IN3(n1938), .IN4(
        MulCntrl_Debug[3]), .OUT(n1937) );
  AOI22 U2013 ( .IN1(n1939), .IN2(AdderCntrl_Debug[4]), .IN3(n1938), .IN4(
        MulCntrl_Debug[4]), .OUT(n1940) );
  NOR2X1 U2014 ( .IN1(n584), .IN2(n1941), .OUT(n1974) );
  NOR2X1 U2015 ( .IN1(n587), .IN2(n2061), .OUT(n1971) );
  AOI22 U2016 ( .IN1(n1820), .IN2(MultResult_reg[0]), .IN3(AdderResult_reg[0]), 
        .IN4(n1821), .OUT(n1942) );
  AOI22 U2017 ( .IN1(n1820), .IN2(MultResult_reg[10]), .IN3(
        AdderResult_reg[10]), .IN4(n1821), .OUT(n1943) );
  AOI22 U2018 ( .IN1(n1820), .IN2(MultResult_reg[11]), .IN3(
        AdderResult_reg[11]), .IN4(n1821), .OUT(n1944) );
  AOI22 U2019 ( .IN1(n1820), .IN2(MultResult_reg[12]), .IN3(
        AdderResult_reg[12]), .IN4(n1821), .OUT(n1945) );
  AOI22 U2020 ( .IN1(n1820), .IN2(MultResult_reg[13]), .IN3(
        AdderResult_reg[13]), .IN4(n1821), .OUT(n1946) );
  AOI22 U2021 ( .IN1(n1820), .IN2(MultResult_reg[14]), .IN3(
        AdderResult_reg[14]), .IN4(n1821), .OUT(n1947) );
  AOI22 U2022 ( .IN1(n1820), .IN2(MultResult_reg[15]), .IN3(
        AdderResult_reg[15]), .IN4(n1821), .OUT(n1948) );
  AOI22 U2023 ( .IN1(n1820), .IN2(MultResult_reg[1]), .IN3(AdderResult_reg[1]), 
        .IN4(n1821), .OUT(n1949) );
  AOI22 U2024 ( .IN1(n1820), .IN2(MultResult_reg[2]), .IN3(AdderResult_reg[2]), 
        .IN4(n1821), .OUT(n1950) );
  AOI22 U2025 ( .IN1(n1820), .IN2(MultResult_reg[3]), .IN3(AdderResult_reg[3]), 
        .IN4(n1821), .OUT(n1951) );
  AOI22 U2026 ( .IN1(n1820), .IN2(MultResult_reg[4]), .IN3(AdderResult_reg[4]), 
        .IN4(n1821), .OUT(n1952) );
  AOI22 U2027 ( .IN1(n1820), .IN2(MultResult_reg[5]), .IN3(AdderResult_reg[5]), 
        .IN4(n1821), .OUT(n1953) );
  AOI22 U2028 ( .IN1(n1820), .IN2(MultResult_reg[6]), .IN3(AdderResult_reg[6]), 
        .IN4(n1821), .OUT(n1954) );
  AOI22 U2029 ( .IN1(n1820), .IN2(MultResult_reg[7]), .IN3(AdderResult_reg[7]), 
        .IN4(n1821), .OUT(n1955) );
  AOI22 U2030 ( .IN1(n1820), .IN2(MultResult_reg[8]), .IN3(AdderResult_reg[8]), 
        .IN4(n1821), .OUT(n1956) );
  AOI22 U2031 ( .IN1(n1820), .IN2(MultResult_reg[9]), .IN3(AdderResult_reg[9]), 
        .IN4(n1821), .OUT(n1957) );
  NOR2X1 U2032 ( .IN1(n1820), .IN2(n1821), .OUT(n1958) );
  AOI22 U2033 ( .IN1(n1820), .IN2(MultExc_reg[0]), .IN3(AddExc_reg[0]), .IN4(
        n1821), .OUT(n1959) );
  AOI22 U2034 ( .IN1(n1820), .IN2(MultExc_reg[1]), .IN3(AddExc_reg[1]), .IN4(
        n1821), .OUT(n1960) );
  AOI22 U2035 ( .IN1(n1820), .IN2(MultExc_reg[2]), .IN3(AddExc_reg[2]), .IN4(
        n1821), .OUT(n1961) );
  NAND3X1 U2036 ( .IN1(getdataStat_reg[1]), .IN2(MBUSY), .IN3(n1767), .OUT(
        n1962) );
  NOR2X1 U2037 ( .IN1(multStateMC[1]), .IN2(n1962), .OUT(MulCntrl_valid) );
  NAND3X1 U2038 ( .IN1(n463), .IN2(n587), .IN3(n1761), .OUT(n1965) );
  OAI21 U2039 ( .IN1(getdataStat_reg[0]), .IN2(n2178), .IN3(n1965), .OUT(n1963) );
  NOR2X1 U2040 ( .IN1(n1833), .IN2(n1963), .OUT(N149) );
  NAND3X1 U2041 ( .IN1(multStateMC[1]), .IN2(n584), .IN3(n1767), .OUT(n1967)
         );
  OAI21 U2042 ( .IN1(getdataStat_reg[1]), .IN2(n2143), .IN3(n1967), .OUT(n1964) );
  NOR2X1 U2043 ( .IN1(n1833), .IN2(n1964), .OUT(N150) );
  OAI21 U2044 ( .IN1(ABUSY), .IN2(n2178), .IN3(n1965), .OUT(n1966) );
  AOI21 U2045 ( .IN1(n1975), .IN2(n1966), .IN3(n1833), .OUT(N151) );
  OAI21 U2046 ( .IN1(MBUSY), .IN2(n2143), .IN3(n1967), .OUT(n1968) );
  AOI21 U2047 ( .IN1(n1976), .IN2(n1968), .IN3(n1833), .OUT(N152) );
  NAND2X1 U2048 ( .IN1(CS), .IN2(AdderCntrl_Dataout_valid), .OUT(n1980) );
  OAI21 U2049 ( .IN1(n1980), .IN2(n1975), .IN3(n587), .OUT(n1969) );
  AOI21 U2050 ( .IN1(DOA), .IN2(n1821), .IN3(n1970), .OUT(N191) );
  NAND2X1 U2051 ( .IN1(CS), .IN2(MulCntrl_Dataout_valid), .OUT(n2062) );
  OAI21 U2052 ( .IN1(n2062), .IN2(n1976), .IN3(n584), .OUT(n1972) );
  AOI21 U2053 ( .IN1(n1820), .IN2(DOA), .IN3(n1973), .OUT(N192) );
  NAND3X1 U2054 ( .IN1(n1834), .IN2(n2237), .IN3(AdderCntrl_Dataout_valid), 
        .OUT(n2236) );
  NAND3X1 U2055 ( .IN1(n1834), .IN2(n2214), .IN3(MulCntrl_Dataout_valid), 
        .OUT(n2213) );
  NAND3X1 U2056 ( .IN1(n806), .IN2(u_Adder_interconnect_stateMC_1_), .IN3(
        Booth_Add_valid), .OUT(n2066) );
  NAND3X1 U2057 ( .IN1(Add_valid), .IN2(n1756), .IN3(n1774), .OUT(n2126) );
  NAND2X1 U2058 ( .IN1(AddSelect), .IN2(n2126), .OUT(n1977) );
  AOI21 U2059 ( .IN1(n2066), .IN2(n1977), .IN3(n1833), .OUT(n1723) );
  AOI21 U2060 ( .IN1(n587), .IN2(n463), .IN3(n1833), .OUT(n1978) );
  NAND2X1 U2061 ( .IN1(n1761), .IN2(n1978), .OUT(n1979) );
  OAI21 U2062 ( .IN1(n2061), .IN2(n2236), .IN3(n1979), .OUT(n1692) );
  AOI21 U2063 ( .IN1(n2237), .IN2(n1980), .IN3(AdderCntrl_valid), .OUT(n1981)
         );
  OAI21 U2064 ( .IN1(n463), .IN2(n462), .IN3(n1981), .OUT(n1982) );
  NOR2X1 U2065 ( .IN1(u_ExcChecker_interconnect_stateMC_0_), .IN2(
        u_ExcChecker_interconnect_stateMC_1_), .OUT(n1995) );
  NAND2X1 U2066 ( .IN1(AdderCntrl_ExcCheck_valid), .IN2(n1772), .OUT(n1983) );
  AOI22 U2067 ( .IN1(u_ExcChecker_interconnect_stateMC_1_), .IN2(n1769), .IN3(
        n1995), .IN4(n1983), .OUT(n1985) );
  NAND2X1 U2068 ( .IN1(MulCntrl_ExcCheck_valid), .IN2(n1834), .OUT(n1984) );
  NAND3X1 U2069 ( .IN1(n1834), .IN2(u_ExcChecker_interconnect_stateMC_0_), 
        .IN3(u_ExcChecker_interconnect_stateMC_1_), .OUT(n1987) );
  OAI21 U2070 ( .IN1(n1985), .IN2(n1984), .IN3(n1987), .OUT(n1661) );
  NAND2X1 U2071 ( .IN1(MulCntrl_ExcCheck_valid), .IN2(
        u_ExcChecker_interconnect_priority_reg), .OUT(n1986) );
  AOI22 U2072 ( .IN1(u_ExcChecker_interconnect_stateMC_0_), .IN2(n1769), .IN3(
        n1995), .IN4(n1986), .OUT(n1989) );
  NAND2X1 U2073 ( .IN1(AdderCntrl_ExcCheck_valid), .IN2(n1834), .OUT(n1988) );
  OAI21 U2074 ( .IN1(n1989), .IN2(n1988), .IN3(n1987), .OUT(n1660) );
  INVX1 U2075 ( .IN(MulCntrl_ExcCheck_valid), .OUT(n1990) );
  AOI22 U2076 ( .IN1(u_ExcChecker_interconnect_priority_reg), .IN2(n1990), 
        .IN3(AdderCntrl_ExcCheck_valid), .IN4(n1772), .OUT(n1992) );
  OAI21 U2077 ( .IN1(u_ExcChecker_interconnect_priority_reg), .IN2(n1995), 
        .IN3(n1834), .OUT(n1991) );
  AOI21 U2078 ( .IN1(n1995), .IN2(n1992), .IN3(n1991), .OUT(n1659) );
  NAND3X1 U2079 ( .IN1(u_ExcChecker_interconnect_stateMC_1_), .IN2(
        MulCntrl_ExcCheck_valid), .IN3(n1773), .OUT(n2068) );
  NAND3X1 U2080 ( .IN1(u_ExcChecker_interconnect_stateMC_0_), .IN2(
        AdderCntrl_ExcCheck_valid), .IN3(n1775), .OUT(n2131) );
  NAND2X1 U2081 ( .IN1(ExcSelect), .IN2(n2131), .OUT(n1993) );
  AOI21 U2082 ( .IN1(n2068), .IN2(n1993), .IN3(n1833), .OUT(n1658) );
  AOI21 U2083 ( .IN1(ExcCheck_valid), .IN2(n1794), .IN3(u_exc_check_StateMC_0_), .OUT(n1994) );
  NOR2X1 U2084 ( .IN1(n1994), .IN2(n1833), .OUT(n1657) );
  NAND3X1 U2085 ( .IN1(n654), .IN2(ExcCheck_valid), .IN3(n1788), .OUT(n1998)
         );
  NOR2X1 U2086 ( .IN1(n1833), .IN2(n1998), .OUT(u_exc_check_N45) );
  NOR2X1 U2087 ( .IN1(n1995), .IN2(n1833), .OUT(n2134) );
  NOR2X1 U2088 ( .IN1(n1833), .IN2(n1769), .OUT(n2132) );
  AOI22 U2089 ( .IN1(n2134), .IN2(MulCntrl_Exc_Ack), .IN3(n1996), .IN4(n2132), 
        .OUT(n1997) );
  NAND3X1 U2090 ( .IN1(MulCntrl_ExcCheck_Datain[10]), .IN2(
        MulCntrl_ExcCheck_Datain[7]), .IN3(ExcSelect), .OUT(n1999) );
  NOR2X1 U2091 ( .IN1(n2000), .IN2(n1999), .OUT(n2009) );
  NAND3X1 U2092 ( .IN1(MulCntrl_ExcCheck_Datain[14]), .IN2(
        MulCntrl_ExcCheck_Datain[8]), .IN3(MulCntrl_ExcCheck_Datain[9]), .OUT(
        n2001) );
  NOR2X1 U2093 ( .IN1(n2002), .IN2(n2001), .OUT(n2008) );
  NOR2X1 U2094 ( .IN1(AdderCntrl_ExcCheck_Datain[13]), .IN2(
        AdderCntrl_ExcCheck_Datain[10]), .OUT(n2003) );
  NAND3X1 U2095 ( .IN1(n2003), .IN2(AdderCntrl_ExcCheck_Datain[8]), .IN3(
        AdderCntrl_ExcCheck_Datain[9]), .OUT(n2004) );
  NOR2X1 U2096 ( .IN1(ExcSelect), .IN2(n2004), .OUT(n2007) );
  NAND3X1 U2097 ( .IN1(AdderCntrl_ExcCheck_Datain[11]), .IN2(
        AdderCntrl_ExcCheck_Datain[12]), .IN3(AdderCntrl_ExcCheck_Datain[14]), 
        .OUT(n2005) );
  NOR2X1 U2098 ( .IN1(AdderCntrl_ExcCheck_Datain[7]), .IN2(n2005), .OUT(n2006)
         );
  AOI22 U2099 ( .IN1(n2009), .IN2(n2008), .IN3(n2007), .IN4(n2006), .OUT(n2138) );
  NOR2X1 U2100 ( .IN1(AdderCntrl_ExcCheck_Datain[3]), .IN2(
        AdderCntrl_ExcCheck_Datain[4]), .OUT(n2011) );
  NOR2X1 U2101 ( .IN1(AdderCntrl_ExcCheck_Datain[2]), .IN2(
        AdderCntrl_ExcCheck_Datain[0]), .OUT(n2010) );
  NOR2X1 U2102 ( .IN1(AdderCntrl_ExcCheck_Datain[1]), .IN2(n2012), .OUT(n2014)
         );
  NOR2X1 U2103 ( .IN1(AdderCntrl_ExcCheck_Datain[5]), .IN2(
        AdderCntrl_ExcCheck_Datain[6]), .OUT(n2013) );
  NAND3X1 U2104 ( .IN1(n2014), .IN2(n2013), .IN3(n1768), .OUT(n2025) );
  NOR2X1 U2105 ( .IN1(MulCntrl_ExcCheck_Datain[3]), .IN2(
        MulCntrl_ExcCheck_Datain[4]), .OUT(n2016) );
  NOR2X1 U2106 ( .IN1(MulCntrl_ExcCheck_Datain[2]), .IN2(
        MulCntrl_ExcCheck_Datain[0]), .OUT(n2015) );
  NOR2X1 U2107 ( .IN1(MulCntrl_ExcCheck_Datain[1]), .IN2(n2017), .OUT(n2019)
         );
  NOR2X1 U2108 ( .IN1(MulCntrl_ExcCheck_Datain[5]), .IN2(
        MulCntrl_ExcCheck_Datain[6]), .OUT(n2018) );
  NAND3X1 U2109 ( .IN1(n2019), .IN2(n2018), .IN3(ExcSelect), .OUT(n2030) );
  NOR2X1 U2110 ( .IN1(AdderCntrl_ExcCheck_Datain[14]), .IN2(
        AdderCntrl_ExcCheck_Datain[9]), .OUT(n2034) );
  NOR2X1 U2111 ( .IN1(AdderCntrl_ExcCheck_Datain[12]), .IN2(n2020), .OUT(n2023) );
  NOR2X1 U2112 ( .IN1(AdderCntrl_ExcCheck_Datain[11]), .IN2(n1731), .OUT(n2022) );
  NOR2X1 U2113 ( .IN1(AdderCntrl_ExcCheck_Datain[8]), .IN2(n1732), .OUT(n2021)
         );
  NAND3X1 U2114 ( .IN1(n2023), .IN2(n2022), .IN3(n2021), .OUT(n2024) );
  NOR2X1 U2115 ( .IN1(n2025), .IN2(n2024), .OUT(n2033) );
  NOR2X1 U2116 ( .IN1(MulCntrl_ExcCheck_Datain[9]), .IN2(
        MulCntrl_ExcCheck_Datain[8]), .OUT(n2032) );
  NOR2X1 U2117 ( .IN1(MulCntrl_ExcCheck_Datain[12]), .IN2(
        MulCntrl_ExcCheck_Datain[11]), .OUT(n2028) );
  NOR2X1 U2118 ( .IN1(MulCntrl_ExcCheck_Datain[14]), .IN2(
        MulCntrl_ExcCheck_Datain[13]), .OUT(n2027) );
  NOR2X1 U2119 ( .IN1(MulCntrl_ExcCheck_Datain[7]), .IN2(
        MulCntrl_ExcCheck_Datain[10]), .OUT(n2026) );
  NAND3X1 U2120 ( .IN1(n2028), .IN2(n2027), .IN3(n2026), .OUT(n2029) );
  NOR2X1 U2121 ( .IN1(n2030), .IN2(n2029), .OUT(n2031) );
  AOI22 U2122 ( .IN1(n2034), .IN2(n2033), .IN3(n2032), .IN4(n2031), .OUT(n2136) );
  OAI21 U2123 ( .IN1(n2138), .IN2(n2035), .IN3(n2136), .OUT(n2036) );
  OAI21 U2124 ( .IN1(n2139), .IN2(n1791), .IN3(n2037), .OUT(n1655) );
  OAI21 U2125 ( .IN1(n2139), .IN2(n1778), .IN3(n2037), .OUT(n1654) );
  AOI22 U2126 ( .IN1(u_booth_Q1_reg), .IN2(n1753), .IN3(n713), .IN4(n1763), 
        .OUT(n2053) );
  NOR2X1 U2127 ( .IN1(Booth_Add_ack), .IN2(n1905), .OUT(n2038) );
  NOR2X1 U2128 ( .IN1(u_Adder_interconnect_stateMC_1_), .IN2(n1756), .OUT(
        n2050) );
  NAND2X1 U2129 ( .IN1(Add_valid), .IN2(n1757), .OUT(n2039) );
  AOI22 U2130 ( .IN1(u_Adder_interconnect_stateMC_1_), .IN2(n1770), .IN3(n2050), .IN4(n2039), .OUT(n2041) );
  NAND2X1 U2131 ( .IN1(n1834), .IN2(Booth_Add_valid), .OUT(n2040) );
  NAND3X1 U2132 ( .IN1(n1834), .IN2(u_Adder_interconnect_stateMC_1_), .IN3(
        n1756), .OUT(n2043) );
  OAI21 U2133 ( .IN1(n2041), .IN2(n2040), .IN3(n2043), .OUT(n1622) );
  NAND2X1 U2134 ( .IN1(Booth_Add_valid), .IN2(
        u_Adder_interconnect_priority_reg), .OUT(n2042) );
  AOI22 U2135 ( .IN1(n2050), .IN2(n2042), .IN3(n1756), .IN4(n1770), .OUT(n2045) );
  NAND2X1 U2136 ( .IN1(n1834), .IN2(Add_valid), .OUT(n2044) );
  OAI21 U2137 ( .IN1(n2045), .IN2(n2044), .IN3(n2043), .OUT(n1621) );
  AOI22 U2138 ( .IN1(u_Adder_interconnect_priority_reg), .IN2(n1780), .IN3(
        Add_valid), .IN4(n1757), .OUT(n2047) );
  OAI21 U2139 ( .IN1(u_Adder_interconnect_priority_reg), .IN2(n2050), .IN3(
        n1834), .OUT(n2046) );
  AOI21 U2140 ( .IN1(n2050), .IN2(n2047), .IN3(n2046), .OUT(n1620) );
  NOR2X1 U2141 ( .IN1(n802), .IN2(u_adder_24b_StateMC_1_), .OUT(n2069) );
  NAND2X1 U2142 ( .IN1(n1834), .IN2(n1792), .OUT(n2048) );
  NOR2X1 U2143 ( .IN1(n2069), .IN2(n2048), .OUT(n1589) );
  AOI21 U2144 ( .IN1(u_adder_24b_StateMC_1_), .IN2(n1792), .IN3(n2069), .OUT(
        n2049) );
  NOR2X1 U2145 ( .IN1(n2049), .IN2(n1833), .OUT(n1588) );
  NOR2X1 U2146 ( .IN1(n2050), .IN2(n1833), .OUT(n2127) );
  NOR2X1 U2147 ( .IN1(n1833), .IN2(n1770), .OUT(n2128) );
  AOI22 U2148 ( .IN1(Booth_Add_ack), .IN2(n2127), .IN3(n2051), .IN4(n2128), 
        .OUT(n2052) );
  AOI22 U2149 ( .IN1(n1904), .IN2(n1796), .IN3(n1903), .IN4(Add_dataout[6]), 
        .OUT(n2055) );
  AOI22 U2150 ( .IN1(n1904), .IN2(u_booth_A_reg_7_), .IN3(n1903), .IN4(
        Add_dataout[7]), .OUT(n2057) );
  AOI21 U2151 ( .IN1(n1767), .IN2(n584), .IN3(n1755), .OUT(n2059) );
  OAI21 U2152 ( .IN1(n2061), .IN2(n2213), .IN3(n2060), .OUT(n1513) );
  AOI21 U2153 ( .IN1(n2214), .IN2(n2062), .IN3(MulCntrl_valid), .OUT(n2063) );
  OAI21 U2154 ( .IN1(n1755), .IN2(n1767), .IN3(n2063), .OUT(n2064) );
  NAND2X1 U2155 ( .IN1(n1770), .IN2(n1834), .OUT(n2065) );
  AOI21 U2156 ( .IN1(n2066), .IN2(n2126), .IN3(n2065), .OUT(
        u_Adder_interconnect_N53) );
  NAND2X1 U2157 ( .IN1(n1769), .IN2(n1834), .OUT(n2067) );
  AOI21 U2158 ( .IN1(n2068), .IN2(n2131), .IN3(n2067), .OUT(
        u_ExcChecker_interconnect_N53) );
  NAND3X1 U2159 ( .IN1(RSTn), .IN2(n2069), .IN3(n768), .OUT(n2070) );
  NOR2X1 U2160 ( .IN1(n1793), .IN2(n2101), .OUT(n707) );
  NAND2X1 U2161 ( .IN1(n1754), .IN2(n1762), .OUT(n2094) );
  NOR2X1 U2162 ( .IN1(u_booth_M_reg_2_), .IN2(n2094), .OUT(n2089) );
  NOR2X1 U2163 ( .IN1(n2090), .IN2(u_booth_M_reg_3_), .OUT(n2085) );
  NOR2X1 U2164 ( .IN1(u_booth_M_reg_4_), .IN2(n2086), .OUT(n2081) );
  NOR2X1 U2165 ( .IN1(n2082), .IN2(u_booth_M_reg_5_), .OUT(n2077) );
  NOR2X1 U2166 ( .IN1(u_booth_M_reg_6_), .IN2(n2078), .OUT(n2073) );
  NOR2X1 U2167 ( .IN1(u_booth_Q1_reg), .IN2(n713), .OUT(n2071) );
  AOI21 U2168 ( .IN1(n2073), .IN2(n1771), .IN3(n2076), .OUT(n705) );
  NAND3X1 U2169 ( .IN1(u_booth_Q1_reg), .IN2(n713), .IN3(n2072), .OUT(n2075)
         );
  OAI21 U2170 ( .IN1(n1771), .IN2(n2073), .IN3(n705), .OUT(n2074) );
  OAI21 U2171 ( .IN1(n2075), .IN2(n1771), .IN3(n2074), .OUT(n704) );
  MUX2X1 U2172 ( .IN1(n2078), .IN2(n2077), .S(u_booth_M_reg_6_), .OUT(n2079)
         );
  AOI22 U2173 ( .IN1(u_booth_M_reg_6_), .IN2(n2097), .IN3(n2098), .IN4(n2079), 
        .OUT(n2080) );
  MUX2X1 U2174 ( .IN1(n2082), .IN2(n2081), .S(u_booth_M_reg_5_), .OUT(n2083)
         );
  AOI22 U2175 ( .IN1(u_booth_M_reg_5_), .IN2(n2097), .IN3(n2098), .IN4(n2083), 
        .OUT(n2084) );
  MUX2X1 U2176 ( .IN1(n2086), .IN2(n2085), .S(u_booth_M_reg_4_), .OUT(n2087)
         );
  AOI22 U2177 ( .IN1(u_booth_M_reg_4_), .IN2(n2097), .IN3(n2098), .IN4(n2087), 
        .OUT(n2088) );
  MUX2X1 U2178 ( .IN1(n2090), .IN2(n2089), .S(u_booth_M_reg_3_), .OUT(n2091)
         );
  AOI22 U2179 ( .IN1(u_booth_M_reg_3_), .IN2(n2097), .IN3(n2098), .IN4(n2091), 
        .OUT(n2092) );
  MUX2X1 U2180 ( .IN1(n2094), .IN2(n2093), .S(u_booth_M_reg_2_), .OUT(n2095)
         );
  AOI22 U2181 ( .IN1(u_booth_M_reg_2_), .IN2(n2097), .IN3(n2098), .IN4(n2095), 
        .OUT(n2096) );
  AOI21 U2182 ( .IN1(n2098), .IN2(n1754), .IN3(n2097), .OUT(n2100) );
  NAND2X1 U2183 ( .IN1(n2098), .IN2(u_booth_N258), .OUT(n2099) );
  AOI22 U2184 ( .IN1(u_booth_M_reg_1_), .IN2(n2100), .IN3(n2099), .IN4(n1762), 
        .OUT(n698) );
  NOR2X1 U2185 ( .IN1(n1754), .IN2(n2101), .OUT(n697) );
  NAND2X1 U2186 ( .IN1(u_exc_check_StateMC_0_), .IN2(n1834), .OUT(n2103) );
  OAI21 U2187 ( .IN1(n654), .IN2(n2103), .IN3(n2102), .OUT(n622) );
  AOI22 U2188 ( .IN1(u_booth_M_reg_7_), .IN2(n2113), .IN3(n2112), .IN4(
        Booth_datain1[7]), .OUT(n2105) );
  AOI22 U2189 ( .IN1(u_booth_M_reg_6_), .IN2(n2113), .IN3(n2112), .IN4(
        Booth_datain1[6]), .OUT(n2106) );
  AOI22 U2190 ( .IN1(u_booth_M_reg_5_), .IN2(n2113), .IN3(n2112), .IN4(
        Booth_datain1[5]), .OUT(n2107) );
  AOI22 U2191 ( .IN1(u_booth_M_reg_4_), .IN2(n2113), .IN3(n2112), .IN4(
        Booth_datain1[4]), .OUT(n2108) );
  AOI22 U2192 ( .IN1(u_booth_M_reg_3_), .IN2(n2113), .IN3(n2112), .IN4(
        Booth_datain1[3]), .OUT(n2109) );
  AOI22 U2193 ( .IN1(u_booth_M_reg_2_), .IN2(n2113), .IN3(n2112), .IN4(
        Booth_datain1[2]), .OUT(n2110) );
  AOI22 U2194 ( .IN1(u_booth_M_reg_1_), .IN2(n2113), .IN3(n2112), .IN4(
        Booth_datain1[1]), .OUT(n2111) );
  AOI22 U2195 ( .IN1(u_booth_N258), .IN2(n2113), .IN3(n2112), .IN4(
        Booth_datain1[0]), .OUT(n2114) );
  AOI21 U2196 ( .IN1(n768), .IN2(n1777), .IN3(n1833), .OUT(n2124) );
  AOI22 U2197 ( .IN1(Add_dataout[1]), .IN2(n1822), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N123), .OUT(n2115) );
  AOI22 U2198 ( .IN1(Add_dataout[2]), .IN2(n1822), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N124), .OUT(n2116) );
  AOI22 U2199 ( .IN1(Add_dataout[3]), .IN2(n1822), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N125), .OUT(n2117) );
  AOI22 U2200 ( .IN1(Add_dataout[4]), .IN2(n1822), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N126), .OUT(n2118) );
  AOI22 U2201 ( .IN1(Add_dataout[5]), .IN2(n1822), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N127), .OUT(n2119) );
  INVX1 U2202 ( .IN(n2119), .OUT(n601) );
  AOI22 U2203 ( .IN1(Add_dataout[6]), .IN2(n1822), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N128), .OUT(n2120) );
  INVX1 U2204 ( .IN(n2120), .OUT(n600) );
  AOI22 U2205 ( .IN1(Add_dataout[7]), .IN2(n1822), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N129), .OUT(n2121) );
  INVX1 U2206 ( .IN(n2121), .OUT(n599) );
  AOI22 U2207 ( .IN1(Add_dataout[8]), .IN2(n1822), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N130), .OUT(n2122) );
  INVX1 U2208 ( .IN(n2122), .OUT(n598) );
  AOI22 U2209 ( .IN1(u_adder_24b_N52), .IN2(u_adder_24b_N131), .IN3(n1822), 
        .IN4(Add_carryout), .OUT(n2123) );
  AOI22 U2210 ( .IN1(Add_dataout[0]), .IN2(n1822), .IN3(u_adder_24b_N52), 
        .IN4(u_adder_24b_N122), .OUT(n2125) );
  AOI22 U2211 ( .IN1(n2129), .IN2(n2128), .IN3(n2127), .IN4(Add_ack), .OUT(
        n2130) );
  AOI22 U2212 ( .IN1(n2134), .IN2(AdderCntrl_Exc_Ack), .IN3(n2133), .IN4(n2132), .OUT(n2135) );
  OAI21 U2213 ( .IN1(n2138), .IN2(n2137), .IN3(n2136), .OUT(n2141) );
  AOI22 U2214 ( .IN1(u_exc_check_N45), .IN2(n2141), .IN3(n2140), .IN4(
        ExcCheck_value[2]), .OUT(n2142) );
  NOR2X1 U2215 ( .IN1(n2143), .IN2(n1833), .OUT(n2176) );
  NOR2X1 U2216 ( .IN1(n1827), .IN2(n1833), .OUT(n2175) );
  AOI22 U2217 ( .IN1(DIN2[0]), .IN2(n1825), .IN3(n1827), .IN4(MulCntrl_Op2[0]), 
        .OUT(n2144) );
  AOI22 U2218 ( .IN1(n1827), .IN2(MulCntrl_Op2[1]), .IN3(n1825), .IN4(DIN2[1]), 
        .OUT(n2145) );
  AOI22 U2219 ( .IN1(n2176), .IN2(MulCntrl_Op2[2]), .IN3(n1825), .IN4(DIN2[2]), 
        .OUT(n2146) );
  AOI22 U2220 ( .IN1(n2176), .IN2(MulCntrl_Op2[3]), .IN3(n1825), .IN4(DIN2[3]), 
        .OUT(n2147) );
  AOI22 U2221 ( .IN1(n2176), .IN2(MulCntrl_Op2[4]), .IN3(n1825), .IN4(DIN2[4]), 
        .OUT(n2148) );
  AOI22 U2222 ( .IN1(n1827), .IN2(MulCntrl_Op2[5]), .IN3(n1825), .IN4(DIN2[5]), 
        .OUT(n2149) );
  AOI22 U2223 ( .IN1(n1827), .IN2(MulCntrl_Op2[6]), .IN3(n1825), .IN4(DIN2[6]), 
        .OUT(n2150) );
  AOI22 U2224 ( .IN1(n2176), .IN2(n1818), .IN3(n1825), .IN4(DIN2[7]), .OUT(
        n2151) );
  AOI22 U2225 ( .IN1(n2176), .IN2(MulCntrl_Op2[8]), .IN3(n1825), .IN4(DIN2[8]), 
        .OUT(n2152) );
  AOI22 U2226 ( .IN1(n2176), .IN2(n1735), .IN3(n1825), .IN4(DIN2[9]), .OUT(
        n2153) );
  AOI22 U2227 ( .IN1(n1827), .IN2(n1734), .IN3(n1825), .IN4(DIN2[10]), .OUT(
        n2154) );
  AOI22 U2228 ( .IN1(n1827), .IN2(n1737), .IN3(n1825), .IN4(DIN2[11]), .OUT(
        n2155) );
  AOI22 U2229 ( .IN1(n2176), .IN2(n1738), .IN3(n1825), .IN4(DIN2[12]), .OUT(
        n2156) );
  AOI22 U2230 ( .IN1(n2176), .IN2(MulCntrl_Op2[13]), .IN3(n2175), .IN4(
        DIN2[13]), .OUT(n2157) );
  AOI22 U2231 ( .IN1(n1827), .IN2(MulCntrl_Op2[14]), .IN3(n1825), .IN4(
        DIN2[14]), .OUT(n2158) );
  AOI22 U2232 ( .IN1(n1827), .IN2(MulCntrl_Op2[15]), .IN3(n1825), .IN4(
        DIN2[15]), .OUT(n2159) );
  AOI22 U2233 ( .IN1(n1827), .IN2(MulCntrl_Op1[0]), .IN3(n2175), .IN4(DIN1[0]), 
        .OUT(n2160) );
  AOI22 U2234 ( .IN1(n1827), .IN2(MulCntrl_Op1[1]), .IN3(n2175), .IN4(DIN1[1]), 
        .OUT(n2161) );
  AOI22 U2235 ( .IN1(n1827), .IN2(MulCntrl_Op1[2]), .IN3(n1825), .IN4(DIN1[2]), 
        .OUT(n2162) );
  AOI22 U2236 ( .IN1(n1827), .IN2(MulCntrl_Op1[3]), .IN3(n1825), .IN4(DIN1[3]), 
        .OUT(n2163) );
  AOI22 U2237 ( .IN1(n1827), .IN2(MulCntrl_Op1[4]), .IN3(n1825), .IN4(DIN1[4]), 
        .OUT(n2164) );
  AOI22 U2238 ( .IN1(n1827), .IN2(MulCntrl_Op1[5]), .IN3(n2175), .IN4(DIN1[5]), 
        .OUT(n2165) );
  AOI22 U2239 ( .IN1(n1827), .IN2(MulCntrl_Op1[6]), .IN3(n2175), .IN4(DIN1[6]), 
        .OUT(n2166) );
  AOI22 U2240 ( .IN1(n1827), .IN2(MulCntrl_Op1[7]), .IN3(n1825), .IN4(DIN1[7]), 
        .OUT(n2167) );
  AOI22 U2241 ( .IN1(n1827), .IN2(MulCntrl_Op1[8]), .IN3(n1825), .IN4(DIN1[8]), 
        .OUT(n2168) );
  AOI22 U2242 ( .IN1(n1827), .IN2(MulCntrl_Op1[9]), .IN3(n1825), .IN4(DIN1[9]), 
        .OUT(n2169) );
  AOI22 U2243 ( .IN1(n1827), .IN2(MulCntrl_Op1[10]), .IN3(n1825), .IN4(
        DIN1[10]), .OUT(n2170) );
  AOI22 U2244 ( .IN1(n1827), .IN2(MulCntrl_Op1[11]), .IN3(n1825), .IN4(
        DIN1[11]), .OUT(n2171) );
  AOI22 U2245 ( .IN1(n1827), .IN2(n1817), .IN3(n1825), .IN4(DIN1[12]), .OUT(
        n2172) );
  AOI22 U2246 ( .IN1(n1827), .IN2(n1814), .IN3(n1825), .IN4(DIN1[13]), .OUT(
        n2173) );
  AOI22 U2247 ( .IN1(n1827), .IN2(MulCntrl_Op1[14]), .IN3(n2175), .IN4(
        DIN1[14]), .OUT(n2174) );
  AOI22 U2248 ( .IN1(n1827), .IN2(MulCntrl_Op1[15]), .IN3(n1825), .IN4(
        DIN1[15]), .OUT(n2177) );
  NOR2X1 U2249 ( .IN1(n2178), .IN2(n1833), .OUT(n2210) );
  NOR2X1 U2250 ( .IN1(n1829), .IN2(n1833), .OUT(n2211) );
  AOI22 U2251 ( .IN1(DIN2[0]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op2[0]), .OUT(n2179) );
  AOI22 U2252 ( .IN1(DIN2[1]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op2[1]), .OUT(n2180) );
  AOI22 U2253 ( .IN1(DIN2[2]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op2[2]), .OUT(n2181) );
  AOI22 U2254 ( .IN1(DIN2[3]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op2[3]), .OUT(n2182) );
  AOI22 U2255 ( .IN1(DIN2[4]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op2[4]), .OUT(n2183) );
  AOI22 U2256 ( .IN1(DIN2[5]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op2[5]), .OUT(n2184) );
  AOI22 U2257 ( .IN1(DIN2[6]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op2[6]), .OUT(n2185) );
  AOI22 U2258 ( .IN1(DIN2[7]), .IN2(n1831), .IN3(n1829), .IN4(n1815), .OUT(
        n2186) );
  AOI22 U2259 ( .IN1(DIN2[8]), .IN2(n1831), .IN3(n1829), .IN4(n1809), .OUT(
        n2187) );
  AOI22 U2260 ( .IN1(DIN2[9]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op2[9]), .OUT(n2188) );
  AOI22 U2261 ( .IN1(DIN2[10]), .IN2(n1831), .IN3(n2210), .IN4(n1740), .OUT(
        n2189) );
  AOI22 U2262 ( .IN1(DIN2[11]), .IN2(n1831), .IN3(n1829), .IN4(n1739), .OUT(
        n2190) );
  AOI22 U2263 ( .IN1(DIN2[12]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op2[12]), .OUT(n2191) );
  AOI22 U2264 ( .IN1(DIN2[13]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op2[13]), .OUT(n2192) );
  AOI22 U2265 ( .IN1(DIN2[14]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op2[14]), .OUT(n2193) );
  AOI22 U2266 ( .IN1(DIN2[15]), .IN2(n2211), .IN3(n1829), .IN4(
        AdderCntrl_Op2[15]), .OUT(n2194) );
  AOI22 U2267 ( .IN1(DIN1[0]), .IN2(n2211), .IN3(n1829), .IN4(
        AdderCntrl_Op1[0]), .OUT(n2195) );
  AOI22 U2268 ( .IN1(DIN1[1]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op1[1]), .OUT(n2196) );
  AOI22 U2269 ( .IN1(DIN1[2]), .IN2(n2211), .IN3(n1829), .IN4(
        AdderCntrl_Op1[2]), .OUT(n2197) );
  AOI22 U2270 ( .IN1(DIN1[3]), .IN2(n2211), .IN3(n1829), .IN4(
        AdderCntrl_Op1[3]), .OUT(n2198) );
  AOI22 U2271 ( .IN1(DIN1[4]), .IN2(n2211), .IN3(n1829), .IN4(
        AdderCntrl_Op1[4]), .OUT(n2199) );
  AOI22 U2272 ( .IN1(DIN1[5]), .IN2(n1831), .IN3(n2210), .IN4(
        AdderCntrl_Op1[5]), .OUT(n2200) );
  AOI22 U2273 ( .IN1(DIN1[6]), .IN2(n2211), .IN3(n1829), .IN4(
        AdderCntrl_Op1[6]), .OUT(n2201) );
  AOI22 U2274 ( .IN1(DIN1[7]), .IN2(n1831), .IN3(n2210), .IN4(n1808), .OUT(
        n2202) );
  AOI22 U2275 ( .IN1(DIN1[8]), .IN2(n1831), .IN3(n2210), .IN4(n1810), .OUT(
        n2203) );
  AOI22 U2276 ( .IN1(DIN1[9]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op1[9]), .OUT(n2204) );
  AOI22 U2277 ( .IN1(DIN1[10]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op1[10]), .OUT(n2205) );
  AOI22 U2278 ( .IN1(DIN1[11]), .IN2(n1831), .IN3(n2210), .IN4(
        AdderCntrl_Op1[11]), .OUT(n2206) );
  AOI22 U2279 ( .IN1(DIN1[12]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op1[12]), .OUT(n2207) );
  AOI22 U2280 ( .IN1(DIN1[13]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op1[13]), .OUT(n2208) );
  AOI22 U2281 ( .IN1(DIN1[14]), .IN2(n1831), .IN3(n1829), .IN4(
        AdderCntrl_Op1[14]), .OUT(n2209) );
  AOI22 U2282 ( .IN1(DIN1[15]), .IN2(n1831), .IN3(n2210), .IN4(
        AdderCntrl_Op1[15]), .OUT(n2212) );
  AOI21 U2283 ( .IN1(n2214), .IN2(MulCntrl_Dataout_valid), .IN3(n1833), .OUT(
        n2233) );
  AOI22 U2284 ( .IN1(n2234), .IN2(MulCntrl_Dataout[15]), .IN3(n1823), .IN4(
        MultResult_reg[15]), .OUT(n2215) );
  AOI22 U2285 ( .IN1(n2234), .IN2(MulCntrl_Dataout[14]), .IN3(n1823), .IN4(
        MultResult_reg[14]), .OUT(n2216) );
  AOI22 U2286 ( .IN1(n2234), .IN2(MulCntrl_Dataout[13]), .IN3(n1823), .IN4(
        MultResult_reg[13]), .OUT(n2217) );
  AOI22 U2287 ( .IN1(n2234), .IN2(MulCntrl_Dataout[12]), .IN3(n1823), .IN4(
        MultResult_reg[12]), .OUT(n2218) );
  AOI22 U2288 ( .IN1(n2234), .IN2(MulCntrl_Dataout[11]), .IN3(n1823), .IN4(
        MultResult_reg[11]), .OUT(n2219) );
  AOI22 U2289 ( .IN1(n2234), .IN2(MulCntrl_Dataout[10]), .IN3(n1823), .IN4(
        MultResult_reg[10]), .OUT(n2220) );
  AOI22 U2290 ( .IN1(n2234), .IN2(MulCntrl_Dataout[9]), .IN3(n1823), .IN4(
        MultResult_reg[9]), .OUT(n2221) );
  AOI22 U2291 ( .IN1(n2234), .IN2(MulCntrl_Dataout[8]), .IN3(n1823), .IN4(
        MultResult_reg[8]), .OUT(n2222) );
  AOI22 U2292 ( .IN1(n2234), .IN2(MulCntrl_Dataout[7]), .IN3(n1823), .IN4(
        MultResult_reg[7]), .OUT(n2223) );
  AOI22 U2293 ( .IN1(n2234), .IN2(MulCntrl_Dataout[6]), .IN3(n1823), .IN4(
        MultResult_reg[6]), .OUT(n2224) );
  AOI22 U2294 ( .IN1(n2234), .IN2(MulCntrl_Dataout[5]), .IN3(n1823), .IN4(
        MultResult_reg[5]), .OUT(n2225) );
  AOI22 U2295 ( .IN1(n2234), .IN2(MulCntrl_Dataout[4]), .IN3(n1823), .IN4(
        MultResult_reg[4]), .OUT(n2226) );
  AOI22 U2296 ( .IN1(n2234), .IN2(MulCntrl_Dataout[3]), .IN3(n1823), .IN4(
        MultResult_reg[3]), .OUT(n2227) );
  AOI22 U2297 ( .IN1(n2234), .IN2(MulCntrl_Dataout[2]), .IN3(n1823), .IN4(
        MultResult_reg[2]), .OUT(n2228) );
  AOI22 U2298 ( .IN1(n2234), .IN2(MulCntrl_Dataout[1]), .IN3(n1823), .IN4(
        MultResult_reg[1]), .OUT(n2229) );
  AOI22 U2299 ( .IN1(n2234), .IN2(MulCntrl_Dataout[0]), .IN3(n1823), .IN4(
        MultResult_reg[0]), .OUT(n2230) );
  AOI22 U2300 ( .IN1(n2234), .IN2(MulCntrl_Exc[2]), .IN3(n1823), .IN4(
        MultExc_reg[2]), .OUT(n2231) );
  AOI22 U2301 ( .IN1(n2234), .IN2(MulCntrl_Exc[1]), .IN3(n1823), .IN4(
        MultExc_reg[1]), .OUT(n2232) );
  AOI22 U2302 ( .IN1(n2234), .IN2(MulCntrl_Exc[0]), .IN3(n1823), .IN4(
        MultExc_reg[0]), .OUT(n2235) );
  AOI21 U2303 ( .IN1(n2237), .IN2(AdderCntrl_Dataout_valid), .IN3(n1833), 
        .OUT(n2256) );
  AOI22 U2304 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[15]), .IN3(n1824), .IN4(
        AdderResult_reg[15]), .OUT(n2238) );
  AOI22 U2305 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[14]), .IN3(n1824), .IN4(
        AdderResult_reg[14]), .OUT(n2239) );
  AOI22 U2306 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[13]), .IN3(n1824), .IN4(
        AdderResult_reg[13]), .OUT(n2240) );
  AOI22 U2307 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[12]), .IN3(n1824), .IN4(
        AdderResult_reg[12]), .OUT(n2241) );
  AOI22 U2308 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[11]), .IN3(n1824), .IN4(
        AdderResult_reg[11]), .OUT(n2242) );
  AOI22 U2309 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[10]), .IN3(n1824), .IN4(
        AdderResult_reg[10]), .OUT(n2243) );
  AOI22 U2310 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[9]), .IN3(n1824), .IN4(
        AdderResult_reg[9]), .OUT(n2244) );
  AOI22 U2311 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[8]), .IN3(n1824), .IN4(
        AdderResult_reg[8]), .OUT(n2245) );
  AOI22 U2312 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[7]), .IN3(n1824), .IN4(
        AdderResult_reg[7]), .OUT(n2246) );
  AOI22 U2313 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[6]), .IN3(n1824), .IN4(
        AdderResult_reg[6]), .OUT(n2247) );
  AOI22 U2314 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[5]), .IN3(n1824), .IN4(
        AdderResult_reg[5]), .OUT(n2248) );
  AOI22 U2315 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[4]), .IN3(n1824), .IN4(
        AdderResult_reg[4]), .OUT(n2249) );
  AOI22 U2316 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[3]), .IN3(n1824), .IN4(
        AdderResult_reg[3]), .OUT(n2250) );
  AOI22 U2317 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[2]), .IN3(n1824), .IN4(
        AdderResult_reg[2]), .OUT(n2251) );
  AOI22 U2318 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[1]), .IN3(n1824), .IN4(
        AdderResult_reg[1]), .OUT(n2252) );
  AOI22 U2319 ( .IN1(n2257), .IN2(AdderCntrl_Dataout[0]), .IN3(n1824), .IN4(
        AdderResult_reg[0]), .OUT(n2253) );
  AOI22 U2320 ( .IN1(n2257), .IN2(AdderCntrl_Exc[2]), .IN3(n1824), .IN4(
        AddExc_reg[2]), .OUT(n2254) );
  AOI22 U2321 ( .IN1(n2257), .IN2(AdderCntrl_Exc[1]), .IN3(n1824), .IN4(
        AddExc_reg[1]), .OUT(n2255) );
  AOI22 U2322 ( .IN1(n2257), .IN2(AdderCntrl_Exc[0]), .IN3(n1824), .IN4(
        AddExc_reg[0]), .OUT(n2258) );
endmodule

